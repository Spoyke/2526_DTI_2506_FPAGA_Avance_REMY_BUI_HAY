// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
WTVXbR+zb5ANmqeApCNaWmf/S2jy9k09eugdwXov7oAGtvsfoITadjLhaS0Wb77x4Pd1zfyu2naB
XMU5NbAXvQ5mHq4IieJ+BOXn/TbLDI0IiErSBNEpNxxs+/OzFE4m7M7oPDSWPCMurXm/dEFMjYK8
UhNHfuqkGB0kVflfvZqGzeTMOxrc1dX786DpO8YwFhYNZ3Fr2Sfzed09u8leQWXwG16PtnTOGzEH
k6LP/aQBns5CCXrBhdSj5DtkUkIrdHl9gQjEIZlHrM1YDmKbisCx09T5OmWU+bitcIft4yJdVUHZ
UyJilSY2EElGJAQz5ApNjn9do+uj+a8jd1TlBQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 32192)
ohMFiBYkJp4Fs+ApUiIF7B0fB99LC/3X5CWTwYY8Y0A07ZVQP45MQp0Ka5A6U8GMqvMSIdDzOVL3
ETQZduyL5LAHuhbqHTsxu7nJFSdiXGKiuHt3eEcu8KMgqEAhOFYGEV9vreDlyGzxaGQIipQymWSN
xgjlEeDYw+Tr5I8wosq0M2+UzuffsdHT4wHqI7bYvkTfjD8rVPBUYuSYKFakAAgZX0Nc6tV7g0uX
v7F9GGu5vCLNKDEEcC1oJ5poWx+TaJV+x5CJK2kVFimWgZ/UgUhgOYfegG1SMwM2AP63C9qbowzG
ZXP5nrUotcmxSafv0uhQumlpVOZ28PcUXauvKwyVrV1lXF1zC3IZz0fqeGGFkFedmDKuhL67GBDO
YEbi6mEVWNddWohzkQeJruIYI/XhyduOvyWERGN70hvmiH9mNEkS70r4ftNoRD84k4MspQVGGfPt
Tz92q4Fp7kQbY4fcppBQo6Ko+CHn/3ndctf2mXcAfejaT9aDsTK9yWcgxbkN7Esd+lhDBhEowJ3w
wSvmn5QYFujiOSjtGUMtykILIDSa/7PH7Ar8Cd+2VMHonInMMidfERlN1tNMcKPnMeZCpfD6hW8Z
fabA8R7z62V7U5LyxeA2FmWnKsC3lP7gCKgvDOZMKE6Hk8tsG0hN6jXx+JsaXpmyvVDBqZuhifzr
2rtut0ROoADlFxWk5ruYD2ntaiQhZRmxsyLD6sT35NlUlk9UQ1aT5ptrV00XXReRGC9tcb0+lI+M
gkJAEVfibNqR4ZTlVq/YyR2nP0SRrAp40pYg2PNSe1WkbDWu5J4XWKtW6izAd8FSLXX/pXvOyX0T
UyqEbJXas0mLAFkXBPF3ynCNK8PqEsM05W/Av7H3hsHxNeaH4xhEqa8PPZYDmhrs1CjSyD31R7HM
vwT8ZTF7/ZjNBNNMHaoMWP9v/jyXtN397zme484Iri+Ad4fGLhlrNHy3EMLKgKD980LBDXmWfiUh
0g+99phAhVtfqhUMTSV9ZvNVXqL+8FCci/3Ok2cyHyCE3kiMZfv41qp/Qgo7jEZNyW10/XjbuIPe
Mod+rXk5rL8YVj5Oezs/U/0YVvGo7FxXhJrLSSQuV5lt6bFxZa+67dp3BvqtAUxoT0fKjUoe55P5
jkgZ6QFhs+HnpFcNypDEO/Z27AYxuQmDAZLBqUAbMX2xqkEcDW4bepfKULGX7LHKwCiS6uh/dlV0
OthHycvGaTnZk0aLkWw/4QV7A1D4m4B9kGBSrIKn2jF+dG4iDNPZ70RGwGzWOmaL5/EzD+PPCs1Z
7ZaHT3UX61cxoSHdjBLnOH0mrn06I02YAfHB+FfecyTfDeAEdJABJroK4aVf51N9MeT0ygcDT8zA
mKaj6NHRTLmJyJ3Uyoyde0FTIaBbLFIunjAbvQknnPxRC6U1q7KPDsjZytTzaOeOAZ7kV9UfQJyz
ZJfUp9MDz+Qso0t2QgCOvN2HFlYKLK70DIpgXDuU9zdOsEIRZnmyKdZVHjc0v/1fUcEEtpBpbtiO
8n6BM1rw0UWhVBa+2XLZ00qXLMWDZi8/MJ97MugCVQqjDDeNf8oCeANnzZHH1N/BMO2k8cw7OaMQ
IpATtmd9hbYl8YNOQYo4nJIiSOl9V31b9yrIms9Wu8rWrT+wuKd1LxNV7PjOyvAYCwKMFqlZtIGd
ZiIilncVzqDM3hls8JmWgzcU8iMBjoW+C3nzIpDzoqgGB9hvVnyNLza8nvsySweZjZJPctZAz5Im
9XpWkd3Pq18xvBPQZHJ4aXe8+bB7gcbwGUMNUYnhR1YclTxCIH2ClZ37f3Il5bbr3Hz2t6bKXDci
MzCKDsUvV7Cf4Or/I9IIY0pqArKfxCxgequ+xawlYTSH0c11ar9QX7Dn3C9q7RoT7YS7GddXa8Wf
+kwXxb58H1W3PWgROsE4/ahPpNY7r5o5Rkig5AwFIzOlddqggx2IWO+eL8rdafFicX3WXz5NDUKk
eqUG/WMhYkBla/VDixym/splurMrgfqdTfp7jrzQvO+kF0x0G9oO0T39vLivxz/RAaTzP6fU/tZd
hbYhrShv16+9Rohokvs3gqH1TtLQj6MDE2Pqs5FLba+6K9ACLBz+DmEoz4crd7VfEBEenHW8Jtja
ve7l8WRDwF/bYfGZ103BQlaLfmKPeaMC0mxsC2IqeKk8aXTpvDxjhgruQSQhlspkNfGmrcVZHEd6
9DCBHQaqN0PdbpqaeNfgHTjGkRH+ry2abYTysB86BhdTJR9woQ6GD7EDIxuq3OfcT7FyKnhAKtXA
kqDbIbQY/xJvyFEZ7BHuVhWFeVlLPwER7X0PaLub3/3qb3kWEZBiIY+0eSNJ7D7hzFvjOVcJPmUL
BSuPm8vbQa8XPXKRwlzH5PgCejih+QJsSJaHXMzoOaoKttxZG8M/eDuJs9WuyW0f8Gx7C8tOnqv4
y1TXfwxOy8RzdY23PGrZ/UqTgK6Bq9Gw6e+jT6FdNRTtOnwIzGMG2U5gWgrdq6PIJDrPMyoNpt7E
YL1Xzw1ABTB6yZ6BJN3ZWysJSM95XasvYy7wPPeEDgSAd+fTgj8nRzHwcNtTkD2HepuqwBo2LgJC
kw85nm7XCKX1SanArY7Cx9rNJlNDqqE5G6bJMujQYfbS1xRDILbFykON2qJQHoABr2KTIJkMyCyJ
DgMRME9OL7Sci4x4bmdyduc48hticasbb53W79nu90ji0BH9FNhxuaU0cRH22IO8j/BY+wJt6nVW
G+6jT7w5C/i84ffTsAMbdAvn73C4BvVkvjEYUkqVCpUXR311ehtXCHKmpg9z950nfwBwT4LS/vjX
g4zuK7H3Zg2/2UsG6TrYQ64J3xQNPxkP1E5tjhZLS09cIlv/nG3ZJn6IWZZ8tV8n5ZAw3iTPzqfQ
5U7B2oauDyqfSqyd6r6+/d814JyvIlkw60Fxtpfde8L+qmmSaF21p8tlzvPwpASiCZBUUbvohsm5
TY8RLyYip7XZk4WfYPm7GETYnMmnBH91W3W53JtQe77V1GJ8MVdEJS/ybIr0IcarHJ8ODgKtdVbf
NYXsy8Q9o92OHvp2FZx9qgj4S7i4pyk4B/BcY1D+0zebaCjylbQX542uOL9k2M39d2szlROMZ/Cq
NaBfeGl9pJ1YN7wfeUxEtOxdlezs/mK9qCUIV01KRUwgxthAGrWahZC16bMiY7rg3x8LPqKuI+Za
mn9YJK0XnApSOOl6/ThKB6BPpJpHjfR+1e/OV9Yx5QQZKAf2JvqGPZFqyehGocLflHMocMhPje6z
tyMOnYsy0+h8NpaDDPPJc98yIrtXBC1i4+5695WdYKStHlZwN/Ry/SFMb9Y0DRmrlpWOf2GrNy48
RmHQ7JOK+bYfUe7MnMIDHC2ACBZd4U3mVKJYHUTHb436m5XgMnOHEjQp9DnhieJGkoABsLgJEdcP
BF2ye7NgGMG4s9iwtKZDNrXe6DXYQMNIYhS+Uqo8aiaRC/l6M4/4uSUpFfD1AYjoQ95CeH6BVFnc
kO/BI8SSGaAn0O1dtwb0R70VaaTmLaoVN3t3yUVJlHkaNetRZrRC1O0D4Kw+6akhznurJ5Z3IGyJ
Ca8GCAaO8Im7oBAkX7Usa1AZl8dlK3EJRZlLnGGCtH5Peek5igAlg+vw7ippu5Gn5G0IqSxZzGc2
/fhbuMMJ+pAx6lErXxz4f+3zytcOP9vOQKb/qTfBJacYni6M9h7DJm/PuzBN8+n3ExQ5GK5E5Fh0
E/Y4xxZC2R75uTUymr8z2bdVblv/RzTccp+RK/S04avke2ko6ZGvK1c70g3NHSjKmNaMVb+zD1r6
TxKYtT6UpBC6lyfsdfPYMDZMSVaEgXRUJ7VCnDHOhZR+5A1tQApXslYV9wPJ7TbCfX3O7/q3d0dj
/Fo0sJ+z7J8+NcqDj5SzF0bickfs4di5MrWj3v1NB/xd4kjoevwo6R5k7wFTh30I5HVsa98EBavp
ztKPhEDkMgDUZH0BaSbzdGjOTeAFD+XcFYG3QO0uyH8D5ChL3JDxTl/8ByhzjsydAa1vCddNjI2O
4s9P5g6UxUpmkoJu19QJqkVL2y7Ahlv5J7VLpRuUQ9hGm58lnLMHXEmO8t5p4gaVlpKXkJOXUlgf
WqD0sRIDBQCWcjhZPCI6iXDgjKBI6zGUnTBEwq/gTcCtkyUK9Dq9kWaAxQXTxH2hOezL7DICe3fa
jS+QhyUPEiIeRn5EpFhF/WKmZOcyjkKbdINvwtk0mCWfdYR9iuut6+5BlplsXq0JPtXL2ovlsBib
AxzpRUczl9WDGUnibcMCltOkWIoBI8l7712eBZiw+zPIDEnZ9du/yQbNVAMj7hNTjUNIl/xfH7Bm
3HvEQEzlGD2ul2XYu+qhjYReWuH8YWlmjCi1AbW/1DFtJ5Nz98SHhrg5/5uYZF+kPBpBOmvVDsE6
EGtpERzGEstnSMPetCcyyCPGaCamliXLu+2RP7Dw0zbSftzEI+zeTioESHXyLvsp+XKjuPwuw+oG
83nE0GgFkAPWLsTdK3JYI6VkPGLm9Zie638yCDyuJa18dHI3VCe/Sb9IjAD/DSELXdLw2r5T4fco
Nvzhvty3Ly/cOfYxRnDwav4hjkTpMNddaBisEDVOmWDpZixE2aZneu1AFEWnDBeYuzxJAlmYVuQJ
qZ2LaVX5RnKGE1pdvARCXUbVJQBfafWBoQI1/TVZmnUNUiGLP+NwFovt4azfXo1U/eSkAf5kszci
mWnm7V2457nCMrSurutLpnPJvF8+qAHEk2IIWLC63U/dkTypMPluDFBd0cINS1VhDcXGkIZQd6RV
668K2qAHslr+W1bdVYTkJedqOh4aqAVM1ssli8zNpi6E+s60cZcRyYGX3R4Gmz3nOHBDxvDmQAHM
HZpMNrnnOCN7MOBy9bC1/2bM4VZc5vl5Gn9Zme3NbsNU+yV5syrJPzXR9fOI0vwvsREY/MJD5c/U
UjU0sWP1/x269Ypt1lRDUYY3mYMCTZA8RUVJU6/SV1Yv8O3307A+wKUDPTL6wcpUg1bSM5JLK0Aq
ZSop3nk+9jB6wVHuari6A8UkHNcBXOSxXV0QBY5jmN16BU44Px3N1tX0nrHkjMOLYbpQKnMlO2kC
K/pCczrvQMY/ILvbKZ3LgLXOWVLCO96Bgy0v02cS5ZLCcY1iE+NWXiwAXl0DS2K10953jP3mWXWG
qfAs8Z42DL2Fmsa2eUuhlrJvy5ygkvYCdXKVWLWcvBBrYfBfOsiJ8U5+WA8gEmzdPnnZVq2Zv2Hu
vatVGUK5u72ZVUUMFiRJCngJg9vNqysJHXWwEuDGdVV2aGMb9o3A9DjA5nxiwrVI1TWsYknJZwm7
MDIZbgcpM/vVXYRMlqYm7A+9+iGz9B+OZjbss7Q99I3y+lc+KOwNcNbct+pBW6fqLUD/hkMRbyej
5KH+5xVhPwexWaJgcT7sIc3FpOcNEobH89hGpMl1V+Z72Pffg3jCjkUH3/45WLW1KrvfiqYMXNlZ
ovaXXwWpplo6Y08wk0+a6/IQ5pUXtW5E0tT57UoF/1u6s5cV6q4uHqaHJY1YslVVTgABH4bVvUMR
HYHfrZ47Vhch7v3kjsdhfBYNiuyJbqYtRtq3mEo04HeTjo+YJ5PgSuxndu/dXTKrZDGe9a8AyrOe
XpyglGB1XRQ4Q1dfwFzgmifqdKiA6XlnzqbzLmHdjJkZeWNjL4pj072pDdLsLR/mpeHF8FxUjB1t
KmWRicPAWgfbkgKNRl6o5xJOVihua2M1nNDrvtXWyCedrvUGeVZrgR7oUaz6Z4UzJ9AfQ1rx5hxu
ujqTQnknxluNwA8Q2qUcqcUQ/xJL6xF1WScyNuEAHy2NuDzDrUurLLDjdTF62qraATBoej2+TM/Y
nuxAtmFmKeGcSujXQTGQCoLujQNhl+FDWGMzrR4j8rqqsQvIpeDnRCGRjyjnSH+wImJ2JBkERyt0
tMrF2SEG1jDrxOEpEEHlblEWaWrpQASOYiHIr6EPY11JK1/+TBj9t4op4XVGMDZ+3vNwVQ13j8A8
BWewBCPipaN2EbiQokc5i4EWBXuM3qQ7dfNweLfaCBDPAVTND15xKkxeUL917tQAJocBuRfBKy96
Ezf9nuoZTbkpewKjy6YzCygJVdxDmpX4cgKEPB6Fqls46XlCmQ5sGvhgSp6KLQAkUYRpFocE/6q3
cHNq7iCKn/oe5ettOM9eJ2COg3lhDrt5kJEnze7sfIfKkK74c3D832AkxXXFEUT+q8y7yI5iQ9/C
nxXFjAe3f4x6aL1MNpO2dqFwMugi8nn5jw8a2gtynF0kFzNHmochMUI8mJVMBtpTBV+h/+J0pJoB
NvqaR3t4G/t9pIWjrNxLk53InI6/lKbVYvDZR9vtS1mtRjf14fVG/w7DLaeq0ilmr3lQV4sj6vdz
bYicAXUBCT92N0mCkugv1xkDaQDPXCV/Lr+aBa9AFxgJiAcXyNJ9lVnfUZYjm9ev8Fxc+tE8K8mZ
J27+C6SUHroOHB/IoICg2PGJ04lfseQRCkLD8uI80+Vytp76Q7zJDSNZjC6PSIRPaNQedxJoegbc
QJpWOC9ycwwgpwC5PGiZGSm6leBG/uAi9NdoOIf+GeoWGj8JFPCfLGLTSOL37916+lwcxMWRUIO7
x0xZTOyKLxgVYXzJlHftQ6eNLkhBkDch7ccYRoh48CJ8NBnAfVQDykmmsF36YIMcfO5xKSBy5iHH
zOamLoZHxdSPleukGrCPZ3gmVAt5wl3wLpeUGQ+MODegJBF0tT6bGaSEqMYOqlx5J6ynebUGD1GN
4kWnaXljTlt3+kPdiIZU7zBT+IP/HJPtyYXuSxWX3YCqu3xaxczbTf3vrPkrQQYrBwEJfMHQhbNu
CmJ7n/NmQm3eZsex7wUrE2xuy3gZEAR2RVbSJ+N5AkjG8ekOjqm0D4+oPZLwMyTkcl+wijmxpbG1
D73RtIXXjD9B8RjiQdz+ccA7v2xiB4fA9odLGTlkTAZEmuOOvQd4oVu13LN/I9ssvy61sO3HJYE0
Z2MGOJ5W90z2XXJ17DZA19C5FDErsoVH5p+9twuU0/ii+L2XZIknwKJycknUAm8XeaVgoAgzQObO
0hKVscO+Oqz8q6Umq6XLsnNIqeC/QRD14eC+Nxme+rKErM4eKDhKDSmdoR0o3QcYwEGO8fETC/ln
/8YhApMjoEtr5rcOLQ7/66G4wYcMD4pkT9f8FGiur72E51gjYxeJ3wX4K6GMKd1sJgYqMZgZUCCX
oAB9vXKAW8POH/7cbQgVFzBNQ6DzRYOqbVN/SfVgLi/flJ4MjObUiNGtT/vFbco9PElcmjAla74a
KupZhlt/ILmrGRYNwYHw89BufmF2c/8IDoNfzqs9E58v96848rtMBRDVUF/2IflwVvOs+Qh4NlqE
6tnj6N/vdCwNIN2vOa5pS2Rfu5UBGqgGDNO8U9HM0lPA2kny9oUxk6g0CnTLGxU/CgP1+wfmWYFn
N4/x18CUr1ZHZrISmc8I/X9K0qaPtSwIaDL1Na3j6phtciezozsq1Y9pAtIYtkRjOOoCr9rqT7bg
8icmmr+Q99TBEr+Za9VqpQnHzM9qi9vHJ56AeF6j6OVAvioqF6MF/WcZb95DvIns6mNgcxs9BF41
Rt+m0m2Af7d99dVL474NoukF+8W3EBjCvBhIJ6s46F81Ukev95P4inh8yYpCohEXo/a2ljj0p2wL
V4gbReyrJTchhhWqbb1SbOwY1xtw3Ftn9xZ1zLGiUBnxv0ZSqvVQSYXNvA2mXERQkj90bNl/VRzE
0zM0w+Tk2z4/RJiAmBdLbipLturcmAfEWdM3xLNvWq+9Fk1D5npkLnVCu/mqU+fSEz2cgQ3h68fd
nC2rxhEdQiQuRahzuimitZBUlGdrAiUcbR1Poyc/tTiCiWNf+6Eu3QsPjYq060fUFkoWR3Qkxpqm
H53jF5Sof/HregJJcIH0fbAvOPGOBWBklqPPNSf05l2MECCUcaxWTyCdt1zQPmEDICQ9BNMQTUq9
LkXrVjPwWTXJOdOY/T2vjMpwIxRex75mHNk1bCv+OdpOWLPI1FCGzc19JTI/PqaZMYg3R2MxvYtL
95t0Ql3cjWtG645lMd6iptvLHRpZaOWo/zELMJWxNoUBUhClezjx2yLnAtpZZMkh6X+mRDGwHhlj
ZJUoQ/gNxunZW0xL47F1+EgfKOm0PFTOOL72JQwVen2BzJ57dAfilGN/riqx3JrTwa1N7TDOoKFc
O/yNpulGyXl3yYWS8YiVsFDAL+/S6OotswWj813W0uG47ub69RjNE9YzhkxfxLkBQyIxzrMVxmwR
LvCIWScLhuxQhDAkY8oGBnMtrYZpBBjKMZqQTtuatypze+z9X8Wh+FsqPpm56DSUQTMyaoEAYAvu
Yxa1pdQohlqeM2N9inTsx1rZg5e4raK5RKWiJsR+e3PNEloyysI5Mx/Ze1kj/SQT8NobdIlXiH42
a4lbGk1AGFqFyYIgAhG0fL2ldSE+KfGxWcr40nZYZqANW2OIsu5R0OrS7d4Kcs1OM6S8FgkluEJt
Q9qKnVIZhP14tc9SuOVt6g5CDArNGPSTTRvsvtMqviHlKHuHmrn2H5HVzaFUPw+EZ9IMQQ67PHhA
VqXBHs5BY6b+XzaHzS2mQuF8BVJV0XKORkPWbvOzfrRo6ItMNfsmu/0WUx+sDyJxnPzauNw2Cj6f
m1lPR+0+qi1cy8FbTE5jhk4nOyeE8PTgS0c95k3bIs2C2zU7y+81AzuYSvf1lgBWnZ4GF/aJtG+c
T4tPEOs5TKYGFqWFMZ3YaASaXJsskBxnjji99vsnYSPKVf3fpT9/oZ/n6zDGiMv9LcGf4ItVDg56
wIN/BuOxGBhs5UVWGd8iRzqF1NZS2E9zTlarb9axK0hRG6uhx0hDufV4TtrRW9Zy4RCqP80+r0Mn
v8IXSH5ROQfeceklAPjiQrmPOJZPdQVzhvFluTPj/4HxTcGu+dXxRi+ay1UaJlrFTtGZ5CF21Cld
+zVpnaQAdxRswF6Gkr7D+dJIAPxPYlZRFV0BhQLOXoqj1vzWv8cUVTRKgoi1DOJF/2b7y//lhmTZ
NvwOvGD0zlWR60B78aC9S6SOCmo6cgUkam0Yz+DzweNxmBGc/ECHl5VPnkNz5Z5zA8sgazW7ilny
uvdQyoJQTA1OVGxK9woSf6QtwuSNYROjnAg8f8bZAHv2oHPCwBYAXkoxUBhPtvciq00fNWOQ6maT
QATVxzVXJ+eQL5PS8siJShIpAe4Y0BLR368UeEQ3MLGHOpzYUzJ2+UxBTeUTlg8h/MQu2PRWUowP
Qbx64aFAabS93DYAvTixJdF3eBGvpT8KL9NC+IplGlIpGKNAJ0ykAZsFDRbQ1X7Z60jKpULlmRbW
Rbv3/gLSedYmhHnG8hXLlPQulvYWFrdWQUHDwqU1KaTbXwuFMiSrr+wf0FzbUe51T25zyxIbzkao
sJUCUqxg14wzFyUZWIgyFwPB+Owu36C+/TWhu1j5IoXYSLPSyNSk2hLE/LKNLCxcsFO28+iw31Jr
9eFM2EJVzNcTNPKkzQBu4GJ9QxH5sMkJqxv9cUUjvdw+fgT6OkgIDKaJWTHrJgXgf9xAxBCT3qsK
Mh+VvcnzrkEQsd+9ElP30fhQC3J9aM/OHxXV/8ynL0MYaXJgxDkjwu/+lEuylOUVKmNqxx3Bu4m1
OkPaO39S8mw+FCuY9c62tPf1RpLZQpCmpB7bY1JHpcXqrAVmMI2wmrLVbsV2YYwja3EN6DdWR9Wg
RINujaqp9jcAUNrYXYINA/cgM66Q5mr/P6QIuArnLhGVP63wha+u/bFEWa5feDX514rdpiXojsM8
vu0jH4rMogsdsZMnvPoQEkcx/PtqwjVfT30uNLbEkJKZOxbOckQbkzDGy/eR+fmaCmQ8hXEldoeK
Ms9wwKYDzGXaRlOZdrcX2v/oHZXE5n4aGWeCSJnwmDfdJRBxI5UzkTxyznKP/jw2UH6MY6V9H8Rf
iPH7GGlkfdUMMZlfmy/KHkK2tgQ1pPmRxRYVAI+YbriWKMyBdace79q2lfIhTG4t2MSv2O6EbHTM
JSYH36E0AiMOydA0++xiAw0B8KPMhxCA/iKE30rr0VYgcyj1hSDaoTSsGMOki67S/v2Rw7WzM/TG
2yaAn4y0SdMWKSUYIQUMv2rp4fNWXQGgw//emwNt6XX1nUmriNiDQE7+fWkMboeXXR/S9my9J5dZ
r9VvFrE0hcCaP07S7r4udKrDhJrdsyOFfozfIGnkDG+ozHbG3QZN69lkG2mRL9IelBwkj7J79MJe
c1YVUg0zf9/2UIIGkbdwCFXZ72mXJNrHj9ZCUSqKMHE+Wq3VbfG4FrhwoA40SjkAGzF90nHuUokL
LR2Zpc7hRSqLgnM9Uv+e0kFkU5XtmI0Deaax6ZxqRPWy6T+/6IQP6D8WGH8RMaWtvd4hj5BMZfeB
5YXkPgwE4ihv7OHXh8F+gzEVS6FMZ0kKKzrQYijJG5zhXAChcmWfE95zahCnafFDS8ymvzeS8tt/
ial+TBM5dVL1CmLy7bjZtZI6m6+91sqB0ndFhVxTeYWbfzRbPKjOfAq6E0MFen7HchUdvMnZf4U7
wpjZazswpGR9ISfbA3hT1vVVPiOlnVAjY5eV0SrJbHMK/vu1xxamIKXyhS/BET1F+XlbMeHAjRR7
LVfhrHEvj2HAaI+RhZANgaSaRA5MYnAbdN+dqR3bWFGGSv2GhqsOyl5nahFJ9EBEk4wotmaj8OTD
Npht26E4/F8CJI47FRKbXKVcDurtlkN8TNq6NXpL87eSfQKT+cfe5FBU9EenhvSu/f1wiLehTsui
MjoNjV/48j6Eq/9HRq6Shj46RGd6IBs+tXDtq3KBowu6VwPh/4UWTiUMNt4HBQmLQq5b93JoM0nG
dn0fJlW1cKEoDF6D9k+klp3qL6Zohj5+NUEwYUMfpWFKJBP5U5x0hRxf5QFXfCptkHl9Zt5BrUrX
PBjTCHdwdQCg/zvBhSjgh2TD0kiz//UYJlkanYXKRqne/PuNEHsnwmQWD0TYA9Mj45vxB7viRR4L
05HefX4hXomQu/S18VNfbSfJrLquFDd1xFyzwhAXyb+Q6zjK1wgUiwdk2KC0OZbax8I2OaPnROEr
pGkqNPwu7avAPlDitugRUT+Dl5lRbhC/bxxo0g4Q/JPYWhzK4xX2rr9JFGwzq+2fSWggCCXnlZ5I
/iAX/C/OxhypcVHRJKXyQLouhaBpiAn/xKWPkcogqpLK21V+bc4cEOBxxvdAtLoVBqPNuAUCGYma
12YNuM422YqX+6RD05OFmwThl7xDpPEXX5pFbEZ55Y9qsULSdifTedVgzJk9A2JI9dFhnd+C3pma
TmMbmMcJbm0CYfdOhCDugbIb9sgt0G19qQs7TdxIRf0xQw8OpLwhg0uADPv7g1msm8uEOY3wY0Fz
1BVoEKSt03HqIHxR+vE++A+bhbNFaMJM14526Nc/rOk9JrSZYkgqs9mP/1yMSwMS2bzZhRakWtd1
KpbMu/zpnzf3Cl3Y9DfT9ELRAtcqRncDa+ugvzDE6DOC6GuRJfoAvjZpet4JeS//wDW0iobxwDl7
twUNzD9a1fqc7ljDz9zcd8puZdoBomkMa+3X3rzmqqM1fszFvKaaW7E3AO+hQFenj2BVGrxlX4pv
yLy0SkSPoAOXV1k9Mv8eA58wkLLB3t5q+lBOFjPLbx10JgJpnuL7DfVHDRTmaca/olFLCoQJYJhm
iXyUfhSMyYDO/8cQqY5j/no0dTwQ98cDltGiE/e7xTP02F29n0v0Em4tWoZ3toyU+lWU9q6bkLTV
fNy9IqW+Ma1oNXeUVsaDPtdznXF9uopm9o5u3gS7zCIuIGwTwIgl5s/BybIgadxM3d5gXXgWrsXp
4bSZE4Q8/2IGhsVFb7iElHX1k+5SPqHWuJ7OMMQnjC4koAyTI7ZZwmXkxlgn1sAwjS5J6JlvRo5y
swJ1Ng5LiMx7PmvRGVR2kmnvik9uoHYNKKxUG0ENUUuwfnX50B64XMp9N+5VupCl+sdNnl+NAA9j
Qiv6ru6QfsC7Nzkrn2Ga+lIBSZ5LHyT5SexNS/XXHjxi2kGWq2S0ejfjogddrakQH3oPERVCgHWJ
iniHxSewngayPXwK4AIQU/Dfu0eRNV/mp5oJVpoCuJOGjHsEiqKxM5iDtCH77HDTQkeNgR6EeCOM
iTNUwM7LXptVvXTeNZresmRLExvqencf0vcxtvVjG3ztHuOESk58lW11HAycYV2o2SWEkWY3mlwi
PhK3BTi1Y35ZlcRXj8mlqv/y5kBp0S/q97pwxhL+rgIf94lpluQ4GPNBnQg1DT+fmXam5Hu8M8Rx
zYV2b33MAatSQepX7QE+mFNdzwv86fmDTyTIj37JoE5ZhaGWdR67abffwWkYjvudSKTcBGy+L1Du
L9gW/quNjOhyhmsv1c5E3Os9P1URvg4CS9BBsKAVKNIieR33Z7XCQnwiDqDFPgjUKjqR3HWKhxeF
dToYimGH5cYQZMDfD3P58gj+ZLqogCVyNH5yWTNE0Rr3OYty1lRJ/VUAmTy98dZN+j7K5JFjtX1C
pRK7R6G/T5NHi8zdmOBBy6ShJkg1aTZCd2Tx+AFVz9amJ067qbJ6BNLmIRnv8WkNuYB4/iV7OyF/
YH67jMEWWDVlE8bZ131nIy77UEpWwpDprg62vwfwuoHCu/V58RXocHMphVxLhVVLosfYEtFx8Tgo
sUYor+ZDR5bQXuahh820xS9o34GDMoWRRA7v3lSNDYejdZjd+UGpHMwg8ZKgaxHzftfyvG6JUh3c
ocrHRtriHsZpi/pzd8Id+hAB7WLz9TedRI6LSgh1bvyce0iKgNft5Mj0MTueaLgkcd/QPLmypCfx
9tnfO823a1wbbv4bJ7Q7uN3ZgGVUajz+Smym5VebJOgyECM5PA2Ftu6P+ymejwoKkeDN/Sd3pvTx
onECWFfPOC92p4m5jCDfHSSlTHRhQ0n4lv6gglytIQzLnGdd8+W6zwjVjOC+NrDaD/h/LNG98/rc
KpEGS2qSnbSUxHQFWPVAKIRISqRYl8779a/eiX2SPs9vVDcABekpj14rGcMO53lO0wDBdsUZ8Jvt
wg10B6dQD2k7xZetsx5nr5bRJ9QfDa9P7009wbkSe7X+qyxy913ngnqg/IiiX7rrw4i+F4Oef2d/
wEjdop4+ikuvtFbNq9tUQnWKfOuwntwRx4hfFChw2yS1wmDJLz0vbVswBzfjlsBGmV8JQTEnucce
Pkf7moowQQk1U93lBc8Jna5zK8VxUOhjCMxD5cZ9yEk42qM/Dxyml7DAYiQLHDnJXFpo0C4peqTD
vDW1a1iUcbEdOc+3reoFR7hqOIJg5ULieTfnRT/nUkuT/WH+njln7y8XtPzRYrvMjUt6rh0C8Tg3
bBNqdMH3j9s6jXHzuIHM47V432l94OzLF0gIPIW4MotuzAb0sTLilAINqxdoGVTEBVuqfgaMuv2U
uRaxnCnZdA4thBfS0umzMdYFGlhT+ScDOmrP2mkL3X+Q5Qy7tc+Pxuf2SgSlPK10dg1XKFvtiJmz
EmmSYDlRTzoa/2BO+w72utH3wmV0+WyBlzYOnaTKvzCuhH3sMb8WMKLBy+TIzigCKA/3qPa1PQnw
L7vzV2iAs4WkJ8+M3m0GgmUBwFo5ecBEbEVU6/OYbuuyTwceu+5A9HM6OpmqDPVspe0sul9Y4ILm
EWYmLn1Px+wdWxw8HL2QH77FMur9rfOsRZyZbNns31t0+TKVZioh3efHxdBEgnLflakftRRuRurs
Kvn4GJNJhU/OizRZiFiV2/bYF42alXgzt7waOCDkk2Zp5HxRPZd1lNr2gEW4GLouUoXY/398ZB4N
1WFg4YWMpZCRWwoYdh/mUYChx4lSqDBTbO+hKKlsIf5KBq6xbO+cTI4rHBsFzwkIGnXKhSRdSKN+
YGDByKLziEs17DO1hr7qSM01IPvQ6iN+vbKMNZehGkzLIa+l7oQuMRu3WNnL/sLWABA6mmm/6tGE
iElEO2ERMSWhOw61srypxFjaiQB7A6DV2nE4JqXdlOX2kFdHntb1TmFK84SFQ84ZJ2nquycOLqex
Mc2WNM0woQMGcoCw2fNvp6hZV6ODVMly/amuQ5pBabWXCBu4+IE4UZuU3wJVJKNDtELiHMYegRGl
yOQ/lE1Hb3EWAizDAsLQqU3AUDIS9eFv88ZJGNvkHjz0YcMO6kS4kYNVMydu4TzDjvbxIw3O3E+j
1neOY/yGCRQKTgPD8lNNFb1h8ArSU7o5x0C92BFE8Upox4FVh70DfNctaIhfq9RNFR4JG0ZsIx48
kvNUJXLJoNmQfEguzM5cYP58RessI0uAqKdkvaKkELgjcUGSVuSgcax53DZ4fYEM+oZGTTVCEi4S
CgVZg/xeVeZCuWGvCYEak3b49rKmvT9tNbrQ3F25AivBekZGL/Z+DIpBIco66UEW5BB/GGb/AbKL
qAAgFxtU7CFN13zokXMc0lv/9Ha1X9A5zFMDO9m6x6SOrA+eVODDk354RuU9dgGPJq6ahldmSy/Q
ymiLyyazlQ/Fzt6QgwASCmhguIzwK9Ccto/kYUHIYKlB3gaBzgsuH+GEOmFD2ldzIM8Zk3TM2SSO
Ri1RxKlXDijP7RMHtamIuKnfsvf+Bkr6q29t6Je2Rlmr6i7cfBMJ5U2Ctoe8pmgyraJAdOtqqab/
8A9nISV1tEDof4TDA3YWasrjnHDY41+Cb9nnU7Flla7dRKL8ZE+dTDq7zw5Utv4E/62Vr7aA3DHZ
TJReOk4flicDpKoNvhhZa3njePewJU2+nfFu8XhcZPH8VWwviNr4Trl70xyTRdznzMW8USmKE5Ku
WQ5xxvHe1V+rxQe18Sy4iXZkDU2jHPNd1luYlH3sqQ8o7mZLOrAL87SXDvsQMzJQR4wsdA3WgT7y
HH9ICa+9YXdh4udqHKp7kKyr6gBuHY4BiPqQsLP263b2ATwcBw9PDJ65IoaAi5ZVS+TecleJLBl0
LfLN/Nq1zIXfvVSzmzgUB376WYMYxTPOzXnFFotGsB+/zO6u6vJja5LvwoXIoEDfu/QmlJkP3njw
o/g+WBPY6Aoaz2WO/MlcFZAOFz2HdyPCAjyNNax2RWhFYnLW3fvsvUUciGr5yVFrs9bd39Vhq50y
QQunDtHSPX4ZnOHoXzjNCAc227AlFV0pcueiLdbgDM5HN/60I2ZQmj+GvGw+SGTCl0z1jfftMxgP
CLJrF4ogkSGy7IRJ8xO29ANtb/JHtCBG6HzNzSDzzs+R+gxeojA8dlbz5yyl6V+BOyz/TCY82A3A
3t7LGolSRGN4952OSWNnkAvRA6c71C/pkSvzfWRFWqGB3U3w4UZy7rEk+a70Gt+FLkEdTr2Mvc8R
+oPFqmqhKx3mZLdZfXyYO+rg1Sl06ikIRor73/rRKQjRB8chFj49J3VLvQ6e2a+VJjWEu4UscX38
KqjCEiS3iBs2iQg8nkkkm+xrfp6jrC5AtIAgSMz1O0mlccyb4VRkuWBvOEO7T/i6whGm41rHgRA9
ddzH6ps/XNYFQprzV9LM267hvqWik9sMytB2olaEBm3zwnIMA7ePRfDqi/TtoaurD9Fyz2KCVfqj
deK1u+y/0Iuefc4gqwvzWHtqJ3uSm/Z1vfN45kRXPHxaSJMGq5OIXyRFcCPeUlFhOSxUVa1Y7g/N
A2dAcGVwv/A3KgTET1yurBSs62FCSor5L46POvgsNUOsl2YNGraz1+Ez891UZGdXpuTLkrNBp0Jw
/i/k+bDAQQBunF2FU/D9lMMo573J/kSHtKT2a2Za+lSlZpcb+JMkl/HTUwfeOk+iVr9oL5JuoTyX
JQNJzCvQ7c4x2pKwbcvwiy45ogP/Tn7Z0XpK0baN75jW4JahfSK53Roy1fckYPIv1SPiIXPkic7B
I3kNsDXsMEac74SWC6USWb5d0t3dhCON8NZ0/6t/Kj1mBJk9ZYEdS+CxLBejc7MvV4Rfc9khOz4J
JFKYjs90uuZxYuOJRTJiCBFtav8hToU/gBAypbqUyD9vYphBaBKg40F42PJsC1pPupHyOr1mtgzr
K5gVsO5q+fzLwOfi5sqieloNmBrQkL9y51ulHhbSgP9QrRkCPSoDLCPG52qAMxNbU4Ci/ujXU1NN
3OUoiiPK6rqzF19fTdbEwv4BYA+UObnJSwWa843nOFSqBAsljcIawcRhJEGAFlpSrXeRVbIYrf36
kPcjzQI7EOyV4xpQ9jVy/NTponfOOYrUcWfEYWVMeKYu5Cg5PufE22Q9w28h+h7xatuyCjVdvLRp
Qs5l4k8hiL+XPr+ryEZmbab/tpBXX21ftOVtNgoJS2JFsL7uNT8bQE3inVJcPfsJ51NfX9d0VKUi
z+cvAyaVf+ykI0gdNIH5ExeI7FJqQt2FM5xFO9qJMSrxj/EeTcBqm4jy415RNf5cgbVcWcGzPAX9
qu5HWe/PLfK+fcBDLIDF717dmdRTZfoSDPXLUubqfF59N2GfcA6Mv5nUp0azbigG/8lC6GeCoUsV
61NqmqdPoJcGJFJ718k8nn5s9U0zEG1ua7TYL/ETCnEI8pndUURCRstkQ33NNLmK2ALt7HoO6uG4
LE4JBgboI/Y/hLQI04FESMMG8l8N9ZgB/TZbvOnZ8iK/gwx7aR9QsCusUe8l3rOmtALOJoOY7Un4
RFnG11xb93C9m8u3/XNLWxhP8KKoDHhkQFJel4YaP0165rVcOIM03mUhJTaqO7bAdoYdCKmA72jH
voKoruMEvl9qnG3BVowpV2ZqU2F9FrrYB+8rHt52FupYQKfN+XidWwpytxsK8jcWoxd/DfoykOGV
XKZdU1x8925eb/Ulh3zahxbFTansUuXRygE0ebbiDL/d9mAgK76bOfeaRqmsW5bGXsWMkUviiUlD
Ly/oSLHdteW+DzkAqlVCe+KRRoZs3F7YXHmZgF6Yzj7BCHvu8yvFRfyre+fXPI8K96wpoHrRkbgX
jQXpXvRUBeKHco3IZNAtOAMtj3l56WGBXChWi0X87RyASc3Nfl4y4RAPQ4aWXl0W/LiLSR9+eAmV
hd2gsyGhFYw0N9Knvs/nfb3kAV0MNFpGtgAfQagI6Q5N9P1uVN9QYJS5jEUGLyhjJ7ApN8yF7RqQ
qu2y7ovAcSHSnYnBF0EGH4pgkWZ+Qn4g4om8vqgXlNu7n85QGGgyef8asaQCyoiFWfbJENOJWr5t
ie6FGtq7E157LuFmFKm5cX5uwt6ipVsIH6APEsuVWua00SBMaC0TmJ0YC7NoYYHJ+JDThhmNo9dL
d4ixwkypp4BitnBvSYxUuAvKIlnOfCrbY5+/A+cxnKp14z9yg8k5RYtyFAmdkhy9qkTLDdDoEGIv
nf4qcpJWqS6wRbGvQsZU7PCupHy4kS2BI9rJI8tolgc+7LmXMavbPsiVEwlPfB9K2q07dBNRdDED
M1fDPRxfuytWDswMgBTYLc72Vos04Nm5UCoIvusPOVPe89T18uclue0Gf3w/IC1i4n3WEFPj2M65
EbS2ULUPZIKqdsK72zi4Z4R1BBilC3oQo9ZOfbznnVEkCWwCl39dR2otOjjATEVN5mrPYLtYyc8O
M0gplKgsjPrgwP0E2VWRWinz5gpM0kzWghBV5MtBRxkxktjhWKe+Ivn2DSjinF3TZTrOFuQPjSpi
DVWvDX5L6tV8BSaPJihWPiSFAVct2O0hJTpr78q7sdTp/qfN5Hb/SZH6fhpDBJ8p6wzMevYcU2Cb
+Id/WuGCITfyEOXn7hh0PnIDJDHjjaOGYothGZT9/4elAMe/NJaGzjSs/owCVhqoyWay6F0Dmpot
Y0EGaXQjHVxY5806Q0SpfILdPrVLF/FT3d9ch+RiadWs6WvMEYgTRlh+3V/EiZG1E/ipABeO/VkY
do8BhgUOUczExz84vh2UF/9kTnj/etYVQ80NgZAcf3oeI9iTdnmjVD8paMC1dGOYWRcKZi7h4Jj4
oYzcXF/p5P9tvyHqeKU5GYzS79APZOVLTLNNG4M3kmuN75x+nImfeJy7mAyWE3hl6qnBe8TcrvWl
w3cFXfMOEI8RgEVYzZEUUFFOzDamP4MgYOAfzua+K3o+FdZQGAMADnE7QDUznp0vQPiCabc8tWkN
Tu0wnJLmcTlnKDPoHgLUc2SR+6cmnHxENEIPt7BvQr7Gy0N9+doRo6EdivsmztSxEmHWyvOeike4
LNEyNeBunRyhzrrYLouQNv0QMd+wsM5fLZuGver3NpeQ8FEqEYk0Y9RbtDS2XGd2xLXIv263rptk
Gp8BZSRj51nRj06AYluO9xcUbnxwEwCAd5CqmXBZRsg0UO8Jk10pXjvr8BtTut2rrUIz+dOS/cUN
wCXfJIjgYeyJlx/1PwZYmY55z++iGc7/3VZ4knwXF1s4lQD2oHrsLVLYHlTu/m0Nlpb/VRVZqWMg
BqOPHGNquXSaIezF310umsfl08bx7XLT9YI8rR5z6GhcldJ7C3tdddmcLkhfU1Qwm6FG8tLfIcmO
VUPSG8ObbfFQw3fxl5qY9UNIB75NiLg9O4nYLQHFFDyRSIaUwwQnxLnH4YQAbpakTILgnydBZj95
HyysvYip1j93ixkkABEyFesNq6wTWIL0rWF+LD9Q9FB7RHMTHZMv1UJA0BXA+muxUVzmDSpz+d3A
SNZtnqcY8g32ihkX2aj6CnJ66jrRuPVeBpLv3Ux0tbrfaB7Fz6B0VujkwKIqi3PBGG+C1p84vwhm
rCDPM4MGqGh4bk0i/yNq+SKvF5gEDK2DxaHF88x6zMRVBsTRaKcZrzQR1LF4CSK8r1WPy/cZe6GR
QWzDS76PKGG+1tXhuFrFOnHy6gZKYKl47/BKI9PCxE3ybI9kYeQT9SsImZa+B3j/rVQY9nX93dv9
eJThA4QrIvEfncko0Ish6UgX4NSPTFfRGeomsuKwkxjmv2JFchrcxiFg2fxyu7PNgJIikmRcO5+N
n+vsWSuTfJulFwEhY2V4J1YMqxydFyv0JtiCWJENo4h7EcVmE+G0dJQ2BUNlBT+keu9MpYIYPLu9
eGN+B/NC7S2rV1m1TRGD7ccLeKrqJRkRi8vFhgryeRd51UgMf2LGdvD7aXJNcR0oyhg+e+2+rkNX
lbBbq/h0xJrhJ+IqBuNKZs51olvsVLf4SDgmnBu3HIXM2Cw57cQnNwjFwVGBVNkAeJDluOmPQzFs
n5+pJzLG5zv76pVpGL0R9sjdR4lTvi3Jxcg6y4f6wQgFVqFbkyyeQL4K5qYZkEMXlm+kwyw7kRCN
j9xrDt8Y+wKHOcCpQ9t+aVUbDWrfyrPEkxUhuk8wyWK8rXge7NmT8CistIyIG65X3rfZlTwFDFs2
d7iZ5gX+wxjdU00PpMMa6S00+KEk3vCQDkwMdmjyGo1mR3Xnva2mHfAn8inqL31CvakfanQ9jB08
FiIeoh3la03D3fGUP6T1APY7ZhH2hnPeN1KBGTwqwBBlgWLmdvpc+c37SOqbkdt2YIhsvaFW/NLW
XLXO+o8SGHf/ovmrwPQt28wYQXHepGJxm6l3jHTIMOKaMKQ1P8ZwEIH3P2d3qHnw6xIJuBRFI8Ws
cBy33ac/+YFCDkTqTVTOcF2IPm+rsypiJpJJHM0CTsBpxoEbUHaDrCtz7jqmg1oM8eck37g4ryAc
7cYfMgPMJE3OpeHeWIiKQQrxqiDhSCpQFSHohb3w2t1O5sXLubOH/pCcl8m4RaxbkWcRXsGReLdz
1HJBpY5LmmfqdUP1Id1/BLeDHOBMCuyYTwDgV6K73oqJlcn8jFORJdHiayXwESOL1fq1NF3ri00y
rsX1f4nTLdfCOiRUiaQ15SvS5ahLm/m94le75qOc5lpD4sMXFvsY48Ko4VkAtqCpcUcgl4NFhQa3
g8zWc71L1Cu13ME59zkqTv7eLf2BFbUXpAZKtSttHUrEFz3ak1XX3ojPIH63iZtX8J8cnvH2HSY9
uRNwse6ew++5bmjOw7blo2JThAlECUjRAvLmiGLTX8suozKkU6FFJBPVi1cEm6DWXdwOyx0pPSZ5
STVhNwyxTRcyIkfujW+IeBwdUGU7OqRCd/D22jnM0IMKvosg5CWfbYztrewAisn6QUCHhptCiFj6
/57jY77MkF4OMsQndvxZLmYZOaIObJatOzrpRIouc6Bm74/oUBrF5Q9GI9pKK9c4lHP9QaEI2SR2
PMJTQwZFGBA9RHWTsvcmo89UUm+clYlkXu0p+H+97cvBnqIutc8PTFrRUSlocm9e4zEtJfWgiqzt
Etc8M40gAu0+068kadJEgYhThBTGOcOz8EzS9i3SlCawbLScmrIFffBCpCzqg+fmEGn3QApKJCR0
O9Z2VLRGqFat3KKdCK4mx7DZzoR+09vDc7QXWpjCFJinb06+DbK5DZ3Ox/pQIsOEag3XB4j9v7ta
uwF+bXrVXTSGcmbBPpBTYKREog8nAex7trNm3qm0CitKN2r/urC1nKeLATmlTcRgMRKzLFYPtPgj
+4tTmGCv3LZF9hdeL1XzX91j5Duu5uxRa5smyoNtN9xLZpMAWxObQYghMpVxiFhBemj4mGUbEEox
I1b1eZluIJMquYIPgp25FugEJ5qKeL2Xe5aBIR8YkHmhHJe0hx6pL0UVq8WXsNkbqrgBOVOZ37uh
A0vvnxDukXAdH1l+RUuQKdSW8Z0FkYYfepenASx592WKaT+PtQZ4AZIic7/a/5wCK4BT2q5m8IJk
LYjnoLY+Sd9FY2ec9wcZ4cleJsnVnm94Z1NZLamkbSoiQwh/EEgf5/7PG786UF4gIa7Zoy6Y55nq
sEdyK2iSgK5XnV38LJJ7veXDgEnGwOa6JtAFANZPmTMkrqUmpkoHINlYOnBWQp/Ci/8MNHgVPzNp
HLac5JjlQHRjpsOlsi5bEpKeppNrSwKmMaLeqznqNcmZXWS9wvBYTTYleVLuu/e3UtSs2YsKX7aV
c3qPE5i44WZMu7hSNiz8NVREz4TG3Z+c5UOnRavSHGxEYtKMyo96hyyx6tB+VWhqkhyaaG46eDMR
pOhgJz+9R4TAnNHJYZpWMYkA6rR46+/HYH4xPtq72W7NLPKfRr19Nczi464Z5pFK4yyfNVvWgev8
F7u/aAxEoLn794ciAHXN15tkWrnlUlQwlMx1/CPwMdTKWp1/6YTkYLGgWkXPrqwabvXKhNQJqxI4
UkyH+B1ulHkOXiCvQXGpyzDFlwK/NBJkfjzoJ2/1p7ogxC3juNsDNcqoSJYecEBq/MZDautirwjN
g/6tEfYNr2P8qwFehln4jyYLmd/YYrgSX2L8cubKU96Nc4ZTSg7aIl+cX2wO1FkmVRCfaYFc7Wlb
nNmdxGoaOwExKAPW5fjnTkdkcfa43hxfnhyITktUlc5qnBqJqbGe2pweMN3j0gjrT3bXWsNnpWmF
pRHG4m9yuOnJbR3t6C6jSPS6coEkD9tWS7pjC9qD7r17CP/ChJlKkBOUHVTeww63D7QrvujuQagL
VXBYlOblW/YMSaCeVdsLPwQptbhZB0qqzWmbb6ZUZ+2xptvLYuELvgc7oHCbOwqofObLupBByXqa
xv2qMMVETdSs3wLHZRiV/5QhMxCPJbpSpFX1jxnjwz0Z4aDMKmzRnOeNKcCVmeTEjV61ihSsRtm+
EVCGKeWG4XwhEHUTMJ9w2fyP12AaZFyRGw4h/9xZ2wAavAGW1D7p01+7WGH9ekALr3GLvvjsPVPH
OJtz3EnRdL6H9Wqh8ZWr+1lBZACtQ1faK+7eBdU3WwniyGGKq7uoCtdiCZ0+rb6tohVe8Rk7Bzjc
8eZPBCZMc3oXnpwpqu2rVms/nz3hfYELt9bni3Hz1agUBsCQzuWyM/P5o9pPNCykHCvWIjdSCDRS
/aD9BGCAs44hXqhhLLn1tlZjAGqeKk82m8aL3thZsJl0HcWQqrmhcAK3TaMmY/ePFFY0bV/V/cEQ
HyEBd/pXUfhN+kvhV5FvA+Z4SmM1WZ9RP8Jlx3OCHKcShY4Qa5Pv1KPjRWfYn+h13lrI1/ZshB6m
eNDQSVrILXBiwxbw8xhO4dZ9Q/L40FF88OkRdA/RAxX0CrChLYio3kPUZdW5zuY8I8a1s2u7CY4R
f+LKofHAwbqT2AxLvB75IU7CkmYfNQlm7VPLMS6QD+rQO79UWVoQbwSx+6uFmtwoO02CKY0K0gLm
AT2KR+zbAz6hWOJsUBmBFgqNfxQ4WXfrQgUWTcd35WtcH+UbNEmmK273QdrUDrqnJL8KYd2hvIS0
v/+MO9IP4jAjeC4qjCAmEWIqomPl02nNDROJ4qQ0DCYjnO7u/njadWpAEOHxUe2frxL4SnYkgHNP
WqEXYzt5LByL7I4PvQ35O0pgyz9A3MoTxs7gCpJEzU6Y5w9YR7mYl08pt0vXirITdgwF/XRbmYBd
rqA58Twof0JJ/eLyAHOaVbyKuywcbXfq0qPB9S+xfkw8l67ihgZnBEAEKt4am5uu3P2+Huy8ABEk
/99Wj7GF7R+4jsRnK2fxXFPBXz//l9vRHhMy3rkNo5S4qxFzrokrxP1bAV9MxDqRwm15XStyEFp3
lH9ARtSpL5qPF2dbOqrwCKF6Run2ZLhOIiVpW718zObDMqJ3O3fxLxrgA/kG87Z3q9T+eT5iL30T
X9PMi8HAkgjbSWSIpvI9XBmkF+Y/cD3HYlDqb2QLZr1qW0D3d6AWTPzAueEVV2VbmrkckiV9dqLS
F+G7+k609SPwMqez0f1UbG3fC8sKCi+pcTvM9cGcgRsKgS/+F5JYcrzmgiMSzIK7hXtSbXelegUA
n9mqK1h/sSP3l3kegSAxEcITjKEXiEkxM8VAO4ydKDtrZ/Vvlh8EE6xuKKsWH9M136LoASg0wUai
//jvvvb/ixdJEQACS1kzlgQ4pHml30G06BD8gkxwfRH6BdnIgs9SccwtNweO3kwhjgcdjd28hGcZ
tdyIWdPG2lPazkvtI8vlmWb7aB37yy3SsjcYugk83QTQUFdzTyxTnzBpuj858yB/hcw9oI5BtZdj
EYjnOiS6OovrWxKV1bgx8WdITEDsRYQwPn4o1Dw6H+mK3QXjjpCuP0+6auKLppgLwspNblW96v6z
KTICJrHmlIoX0HJ/V0PWNwlOEYu63AMiW9VktGMoahfnmvy0oK/ptObWLdn0+2MQW4o2QSnMUNNd
9ZOsITCZcF55sYLzqE0i16sZ96VD+H4NDj5NWkqgLctr4hEMiYHf5opEusBXeT5M+seXezzYkB5d
BwB1qaBnwjilE3GsdVUks+uOcvY7zYdZr6zcUB37yq06JRObT7I2za8tt/F5UvJpt+fyQ69XddSN
eNpVhaZHaAdF/+Geq7VfGRBfC+jl/PnjXIc+TM0uLucDMNtnzT8YrHKUY7EBdzjGvIe/wYH0JPn8
2VOQyE1xp3eaDHVIzq/sfsmuF1ozsczzbnJvSQ+eNt+5T7UoVsCtUY6ft0fTzdFvbm176n5ds3R9
ll41v5WVe5ISCRRQv7ctq9frUYnY+48OTJZYnOUHoiQdPQS+uypyP7vm4uaw1kNeQYgfBrGxkBjB
kPqe8MhnlTqRIqMSxupqrpnfZrPpR6tCOtbWrAEDgt+ob4vq2yy6cN9p84JSkntiKKXzXTPX4RNK
l1wdns5W9ANXkLOMeJ2st5kJ051scmkbp+HL0cQiBEwQAEPRxXuUxQGUcZjrUt4XgZK0muOQO9fC
UFXT7F+nqCZJodUbZ6kJjrITbCnug5H8ZGU89QpfHHOYs+s3keWMKK3dWuedkD/MhjBC/dtbTS4Z
C/Pj9NI4kXjhSBtDJHWxjm6Wn7mMkuF2+SKXTsb0dhdCK1yRK025L7KH9c0MEe40ldJTKYUU3xfK
woNs6E3WWAoqWbyyeiXH5TL/iGD+SIXFkx4bTnQs3r66vEzWpS8VB4DtavOfoHGNv08qPyn2QD+B
JpFQfTidJ8NDwrg5H7QjPeliXLh11LxBIYLeW8itsw/EC4xpvnkoEWhckI+vvJB/4G1WlLeo2Cnr
Xz/xMMb35SkslCzpJzKFJKv6BFX4DBkJd9NyamVadKjUD0inxHjQUbNSGfc6IZz00Bex5Htp7f5d
3oN4OpGWQVv9oxU/+9Ty3R7au52kgAX3fy7opyqpeS/wNxX8utOOL8CfMTPjj/zQcLAnsv0rKw62
S26YahZQNc/CUrzEMhweebziozFdsbvkz/FkKzhWXAQQdviJYZFixHb0Z2Oo0Izye//0s0ktLNUw
2ccY4jznXlbKHehzjDKDnH68ePOLdjruL6jxctvsG31Xr4FJm65vdEtRu8E76EbExYu/TegwMVQt
kOsTpMqfRy904B3gdhV3uNCACEzSI3iBhNuUnxhywhz5VZohDR/ntw7ItUycsOpGodePMHa1Zhp1
8+SPnjH2tpJh6ajLU+zNaq2n3O59j6KcCsc3hPO85cquQ406L8bmj7CVaxpjDgcJ8MorejYYFawa
bZkPgwwDJHJ9jI9eqj1AX3pCSQufz53+Q3hXWJtbS03IHOEujNLn5DarsKWk486Nt6+acj098Zrf
f9ocpIrrK+YmbcjUOzoVbbo8kqiVcIsKyZl33qYhC2nnzv6wc6xQuJyLqF+BEReSO+Xqb7rIpQYM
VQXLYfgstLrrSF/OstmQRZCHU9APFhZk0vZlNtoPfLeU9PFjMyZ8YvtxmUR/u+dbOH0A12I9+DmZ
69OeyMb6F0kwSMLkGI2dJcso30nVni1rUzRUENrVpNm7vcH7PUmDbbls16i+1zivSA/l+flQilin
qfuMJfRpa8DbdR9w50BzlkARq8OWwew11E/s8FKcNG+sJDnlqrNKWtAou48U8vSNeRjaBvm3e94L
EaP+gXV3s/pRVAuZBdIRjg/mDe9mCj04eQrngftASv8f66EO/FuMwUosSOp95V8kGEf1FA67wP4q
Ro5iZdx/zW7A8volO4WdMvw9HHXdzURwEU2YmbSYmTnSuzjY+GdYf4Uw7ea/x/tbQ8omYWlrpCXx
a39xYkcFbPTHIQvFtEgAqc5bNd4Kd1USHqdZLDKmiPCbJkaqHVhuZ2j4X7E6bKt/74gUY7HtXbTs
mYbQZjOReqnx1TumKshzmDM4hHeTBc8JcHWk15bgD/3FVpuwFmyu3l5NlTfyzOcmxryuqTqaC4ZI
wjPRC1biM4JMghgSp1oxAlCgMsPmGF1G05dkQbB2EnRbgEB3JfbTOCf3mcVkEtq1xTmNWwfKe7Na
jqj6n7gMYbadcDQUyf5I6Xny7hlSPuf2E226nPK8u+mGxv7SC+9oJoj5XBMdMJPsenHCRi8JEV66
cxqOIfOQZ2p0GZRNTaFKcQT3JEu+lBht251dbUet006ZktbzDnOKGy0wHYieiEVL3pNuZotRvKGE
tyTHWXa250htYO52TI0hMCt1ORw+G7rgheu79g0HOmQp170tUxlolzkH61lvnBUXmUKOnknumrUm
Oh+KbIEpSIjvnoFsivji5fxwxtx/kr3JN8d/fqNhPnzq2d51f7B3RHes8IoZAgT3ZPTN/TO+9Yfc
Er0myByCkLvfBSe46CJ/hMiFUhtZxbq0iBxsauJak5BcYch8Uah0blMD+ZTL5p8/+HFMef67GDNR
+unbWw/yIekSOZGO2PwPssuzdeFKTuAJlkP4XgrWm8mVuzkdGXD3OdxLZffD0sQalEn/8zAjY/Tu
SR4PfbIzDnNR4KAsLjulkKafTMU/lh+Ai0ia7ZdV5hVYb/XZ6N+1crcFIAgf+aBDO7D+Vf2jzv9K
dCGUk6z4VvERUUX0jMKTF1mg9lFmNdbMOcItTNcrFtPN3Mo4NDMi0bMFHDfYqZ/nEufXGvpwzSdX
J5AKrDZtqMVcORTUqraRtX43Le6qJe4mTBQjgDZhaNrx0OofiUi4MOxDOP/rql/uGnZI3lNfzEan
/8YYzM8RKLCoAVw4eXP7rTb+wcYgvTt91XUkbq2iw3k/srNHG1onteQmW6S0Md3vbCt4pJkcUsLT
933XbAIOBeY8xyoMkvTUE4PfbNq9LolshnAmj+KgBQImdYlHGx8Na3lUGWvEb01/Ik6QQIKGJb26
zHvC10oeCFuzC038BLiN1oLmiLv2jHW3jEXNf1bX2UX07AzZ89RRD88kfKtweJIol95sevX8auZR
VRO+UT6EmupCrtw6BvMY2hLPtGIY6px8kitwLC2jmqcYhazoYQEdtkKS3w6+duqM3ObN7Ewa2Mb5
jSnVJgp4Wr1WY7gRL2QxY1gidmX1KZQ3JlOtN2cNO6SRixxqFJmzZIxgXsF3Af+PRMu3t/swM+zJ
Rxb9cfWRxrHB4V5/LG4wryDSGWEoIFlGwlB2ZZG92PE8BsQmJUagZ2yFbOVowGU/GgGTPKOdI+Df
FqfBLpgQyiiUOAqFHrNSipcwCd7CUde3ajwpQnwz375e8AH9Ad83TyWNd09G3Wp3tu1QuRitteFm
PaBGFBGfLh7Qu1cmrcCDw2HmytSd2rWgeaU78sGEhOnQ+ZPeNqr0A/83a7Hbwr18wZybHb5yKbes
AnC8/Egq8wWeFf0iPaT+2rCxlOmWqPSLINRHEeQUfZPXhFDQj9K4gCHyrjc+PlFGK0vMokA56KI5
mrXZtVKXqzmhpVJDj1+oVGcIUocVkgZop/02QO5F/dOvbbJzd8K/vbcs+zhPGOCzK9z3cpaZDv1n
fQJThK/gktZzOw1qiQV/LZSK4K39BuogHngLGWhSSItBYzDf1KXPU/Dq52dyU1SVzaPB7GoboKn9
6VFAm5fxDZb6/IV8A69FtnU0VEZfvSDuWfdESXVagg4VUPeK2sV6X8ZAjLvmnYzkLVtQnydcy5yz
grlY9hl8qZm38vVJQYJMYE61XjMAfjhevZ3B74o6LMe4vw1v67W+GsUfJ+1uJrebGx57F/YsXq28
cAe6GcZcJoV78nLmEK2y4CJ5Tr4xYk+RohKvva8EHcAWFWS63ERiHtUzAL+A8sbY2OjFIYBIK6QT
0+ZTI1yWrz3WJhqcuP8+tGYwTKzJHExhc5RhmZ/Cn6223sSxFYMZxIPXzZYhqTSHJjdEsYK7wkyk
q8gNIrenWP+paQYc/hPMamr+80o4KLUB11uI4Si6zKrQsdTofY9BCG2BIajHM9rpp2WFCMPFUFVm
A/dAb5DvQfM/UDhTFsMwduT3c5UW4uIirDsUVcFhoxwJJqJb+oCxhkketANfxq02Es0mdmP1eW6Z
gAdbVthoezbne4uRB9Y8gljcjhf4AENQbkXDTX+I0Q792cchHYuSBkrKuVnEh/kkTY4V0sc7em9y
Fg/EkKWLULce+ZDXGee/XcMWvuORIqt7j4u9uBRlmm1+J7yaRTh+RiBUXDwzHN9Khm6mobn9XMOJ
JB7M2seFQC+yj3QElP3XQvvZQm3pu81+oqygrgMNWISbcYU8gty0bJjJ7i0bhVJJxjM+FN1lujAF
dNDJDnn7HnsyX20s008Y2b8s21TO/avimvWMpbqQy5rGgMfn2csjGHAF7Zc4DyoneU5NYNqn55LN
kw0KEmimubuBSyB00xAzgITrg+wUAyz13I4inHUOn1nvVIr27aSEnG+8TN2o0jGp9EzuUxBg2eRG
Rs5Hrp1KZRBgui0GiO84yVuiCUN8a7zQcqowgaQVUEPMTLs3HdKkODxUpO1MPVt4fPeeqKQ9UaAr
0xplOcq6zja3IEM2y9KDwj0kTksdRmxHUjqP8sd24IwJQBnXjKlKpHomBpoGMi0GE6VAoe8DXPbX
/PGsCbmI++khI8Th46VsoUfkZoFT/C9qrTtEXs/VPHmBtFtQf7vy1B10Iu1yl+GFoWPnFY8x8/N3
5Sl7Lxax6Mg2B2ACyh+OfleQ1QEsKc6KNzFK1EmGc+aLWBCtotszW8P7r8QmKRvjfqJo2sjb6Wxq
YCt9JwYjjnt4jhBKark4/Axv2EZk3Vu8JgAU3eZIAs/dds+AASwDcbKNrjKvUD6gskAu4kAW/2ok
uAJg8WGMmecspeI+DQLXHTG490+M+TruKTgnMmT14hJ4jpns0+qxy4IoR9TzZKsKSkIX493n1/GF
F5QNjMJkXKR68+uOHOcFMFLmH+GiN/d4Uiiv2rrstoSU77Is3/QFm3pUTQnJet9GRc6JGz6fUqg8
xAGIdZddKoHarvAz54qA6v0aIPYxhUUp2AyaluBQyOQE3ooyrW+3p94Luu59bdhvfUeI+VKDjRar
PGczpSc7fU2pr7fhMwZ0x9a7gSt4QRwyQtI/BU00htSaIiGOo/FCPJtdP+UsMgSR98tuiYteTI+j
APy+Sqno4LEuAefb3K0vNGHjnma0Gpj/cF05TSnpmrJR3pLf/b1BOZDIBUfdLnkWW9sm7+vkQLiC
vso9BHP0ktvFckWdhhDvrFgjQhfOzLXPFvKbLfktZKJNawPtAhuqKrn12SjQvKeytRdH2rfSGVal
ZaQ9H5L5FwFK06yMeTOnAo2IoqWm62f0vVFn5Krd9yLoR8i6lGmzke6zmi2L5Um3zTwJh4Ta6Iju
IrQ4hunOtV0Bgk7iq0bw1OAnkIg3HnLj93Ppwc1TGkO6XmOV1JHC8bHalBkG9ZzWw7eb590QgiF/
xbQfsO+gOHW2p2je4xlqXdbhKnfUWhwRAIMLslINHU1nD4PLlcU8agYChhoi2FYmrHv5CL3oNE48
Yfcs64PywF6f82Nn9Vol9cdmBXJhyR6TAFxGz6HjA8vfHjDOiyEErcbtFhX+pJbyB9EoMI4ctkoe
8OVMbGpc3D28XNJClPyHbXH7RWl+YlOdYxVRc7nts+pVKnUKLUlZGKDIAbGryZ1r/6GEAnEQms4M
s2MWS/W4mSkpIEwRY79mLu72AgqowHbUidoEKWt6jlRcx+SMsxjeLNQ9LpFMgZohpClTj4pI2O+u
7sgtVI4O8uLITDV48iqgU31JAZ4h7iJ7IF96rTIbg+lr5M/BpGWKqF7mb8iNMboIha/ufbrZkk9t
Jgui2W3Yb4OsM0Ayvjt4VEA/moh4H+N39HVcPh1ZsPIhSAT2R73Unlhe5GCzm/hDAzsRq5wlW9mJ
k6xJhRWyqFl+VSf8c/mOYX5C1WW5BpQT+FozEWJ0r2Sjjsl/+8YOJ/v5AZllwc8j8ErMiuK9Qm/k
5bu+R2VDwamsSRoxfzKA+OpG83pr0bKRDmMu8uhf2chLihNTW98BEhB4bUDLvZAB8NvDp4HaD5Qr
nduxXFuZUgkhZ/A85dnqcSm9UsTFDKWq0btVlQNww+jf6C7up2e+HntXKWijCoA6qAL4r4ZBxlQd
StGqUPKmw9YtdNo8nse/9N/GuFSSSqgXH0lvZwx/XIHGARmDEUn8hejcYSqPK/bZlRHYeFmspau7
HoRJJaRXGRT8UnAveRw8DFZ64Osa6wPjXctFj+/GdMeaz93zqZIxs+DDX4TWt2c+qWCNilMXZ8p0
ML2fxJV5f85cN1KGvEBgT6Yyx7IbH/B0FLvOtXCmg7LQrc0snghBJlMUXvcH/ZJoJJ4dFqe6FlLl
r3yX0QoQydtMKJZRB8ADMAx90txpX7x39rQqkJP7oVtJn5NWxIhnLIp0G9C69aqExU2vNcbo3/S8
cEZwJPHiEpfzapwjjpeNBg9VgWsEmYyM4OgP3NqQcPxaRpTMTZ7lk1PHpUTMdTJo9EHtGjLPGGhG
EfYM1W2muMq2/GhxYjHtenmJuIoXqlmfFKrkei/5pfdjUIxUf4e2Hb1JQcZnKPyOYJHd4Sa/wqzn
GajUvllSHS15e1n9PEYCDlOXsWxb8aYabpNq1Wex29G6m2WnvCJg/Yz9U6/nLhIn4MsrkW2YIB/E
tYYjoA9I6re3vhOJNCJNFjOwnj+fBySdPfHfCrb4uwIZ3i7peNvhhwk3hhjPIEiOFzUK5TtpuMvY
lTcCrMxWQ14mBzCZsPtilqOSGVtGDwSSkFfXEgbs6uyuZLa5BmpLTAiET/Ld9GRTw6J8WkgqGv2q
IKszkh3COquzW1Zcx1/ygejZy+BVA0/ZMRk9TuR1YSOoLd62Z5ez+ZThxonrFQfxA6McNuxeSDL2
b9ZISyKvWYyTCZB1JNJkhz2snq+i6uTzKR0vlCn1tQqtYJsM9xxB5RrV3gRXOWTzWU5xC4/YaUYB
viEdAntM/CgVKA3YAkDmA+MaJqaaqgUO+HzA7ZtPRY5G9ZWDNHgU0bM6YzsUn4bP4pu5N3YahpnR
sbHJzB7sx1qdincpFqwtQMuI+s6eow4m3B38IJL2hJYR9ji6xcFH1Kx3Up2i3Fh4zg8fbFZnaWfD
52H/bi9kcaZ5ncT2fFXE0/vLWQkion2n2kcBUoUR/KSz6dDV5iL2jL2odkPhyKf5ovugEO1s/wSB
8t7pFPHH2ptXHw20ldWa1bZjWO8Qt/vjq2SAk5Axt5W+T4t+8Iujryn13r2fEeG5qQJrFe5SkAlg
ZJhE05G4dhoy0VShYZLrizkF5Wl5u2pqJXdCUo4Wq4sEJJfcf0AsRQuVwveWxqjBidFH/bERFF+a
PFrUkHYacFBcL3Oxt2L/F++9a06JZ+RQHNi3WbQzuMss8gjSyRzC5Khuv261WrfTqINIXbE02P1N
2Z4undW9xF17LL65JuG+fVjtBaMm6H1017eeVUGu94HJwTMAR0rB/dEbzuP5/juo0BaBv3TE5Vkz
Y8k6RvQhQ099hDKtG5n47e0wK1lOyo35dHPuAyVmIR4cdz8QUqr2sclqoDDhhH3rl/xe0gJ0+NlE
tEFe2W1IctSPL9NPCXX1MwAyBSQYxyLIazdsubOP3QFfRSTyly2fWmjhpjSB/hF5fp2AnEGCzxki
pxkRwW6xJI5vcxsMs3tW1lzCqso69968OPf9joywtdR7jRhE9MPTzJRCcslRy6Y3yzFHkBJm/m8j
P4dMAgYrDY6GfrnZr5f5M2Cm4+SEI7FYHZZMkRdwIZEqH40vVky/ej9AjvVIXIDHbh7bW0qOOqoQ
Ke3nItRnXZbe7XELD04FR+z9o0KgzBiKBizDoMZ0FjnOMsPZG+bdnjKs0ESsGfX5M4mzkEl0dbGx
dGajSmuV2rgbrR/SrpMvopjI6/bAZLVn6095rjH2Y22uEZev08mQfLOhha8+cSvrSf0uWnSjdY09
BXsDYIye3xvIXOiVDBisw8jOQGl8QFmgrIAkEsZOnqbAPVbtZOjWB9O3oBY8XXuQy6pM2SuS/ucI
+9pL/8SdgbOFJH6//UG5y363+C2NnBTER70n1RMG30qOcrp+WfqwvUPsc0+RQAcz2IzkSmuq9DlC
ULDjAcNyK42XkQ21vjBLL948L9LLLuVnRZbh4GnQMT9fT1Zs6P+Ie5NU6382+doKEonSrYF/4xFt
mHKFEAzGyGpythrc3SZRreOwWSfzBHoDEiKmAwMGzsmKkC43gE5q/TXdtbfSczlwDkEkU4mY78E4
hzYTWxw901h3GWllHFo08QnYxGK6CWyqhG66rIEfp2EuVt66WP8oIM6QlwAL6lrbxK/ViOr+tfeK
JJadufHX3MUPnHQrhQAaQ72qvknpYtlfoAcS0dkrCOAuctmww8aBfrgZuoefSqeybGcWmFVZ+Nzz
IVrW1GfIDIBHg56uf2jDf5UoFFP2UmJjBUDLvQwv1Vrwq2pdaR8Gav1oXaefI3bP/YcZ7nVb1DH8
qHBuy4ZFqzj6aH2ZiErCAbKU0PjCqdS4RW12scELhF4nhOHogqi0NVIwz0kltu2m7XEfgHWE5mkT
t5vXQ5NX/M76bPaskZtH+Jz/qJXt+JM9p5X0feDsymLmu2a0TaccbMnLv9pR0D+il59HKM3FnwBT
Nf1OPG8529Htd28fhxeFKzp1qP/HVGBRrZ01gM54/qhylZ4hctXAk0IlVeXphEV0VPo6urNTy/fl
BJJQ4VgLITlEEGWk5BUh+gh6tL+pCE+LdPTbI0pxzx9iL92P326kEpNRyix8so97iKZad3knYjQA
N34tiMxC3QJuBVFDtpuiCzeUp7Ybr14WKTnoEeC8UztRhpIjSvcwNdRF5YB5EyQV5Pk5D+8Gt1FG
XFfHysIKYbkpZqWRjpImGc6dH01zK4cXUTQHTeFJuJDS5qIQRx1ee6VlCayakxKu6dfrk2pWqNcI
rHESs/PAWyPmcKRZRu0wG6m1utc9dEbZtxrYN3cXYY34gcj8OzaXa8SfrBPdxHnLIVgEOBleW5HB
+NE596nM+olk/OFIeVf7prp9eipLqS1dFxfY9spbutK6njIP6J1j/9ygHI22ZIgSOR/uDGzr/qYN
NmQuzhxYnMCcvlGVcCFkPk3eHUuXMYxmge1WAPoNy58Es0k3UpXvfoeNCizp5SPwwtgsQnWcW01S
TEvWOrNXPxviJmtpuB/BaF1j7vqMeDG1cQQx+zHDCfj4Mje63cEVzoTdzn1DKv7b9eoersbdGnwy
bHP0r5OmxcsZoYu4pbgBurpE/ZbmLahMUpsx30zeo5y/Z1RJDq3Ah5jXQUe8kIXiO/c86/h57DLu
tCON6HpJBA+cttj0KsIq+zq9l4vzjBXP6+n3MkYe5Vssebu257TuOyMNI40Kdc9DwNzx29GAj41/
i8KBPnay5jj6g/LpjhObd5gzcfhhdmZWKDh87RmjvBQyEajKSIa2clAlglDppqxgfqOcx0+5MQKo
xQdR7va2fZhTf/5OCpc7awzLix6RPeDq/wnba0uBTPNwHOWdIxPhASQsM2477Vb30Bh8XxQg/G46
fBWMlLFo0Fx9JpWePA6GJmU3epadOCtvi4MmpV1bNkH9B79JgqJ2NBJqtYPM8qAkUEEN5HHXDwRN
kPaWnN4x6+QYPDyKUzoFsE5ie9WNjTJ8NV85loldwoWU9AXeugXp9NlxTt/y3ma3TP+usSdMgSEb
7n2VVAOICZCtB5rWy8R/McKed7w/f2tLVOEAyFHzlY9q+LGTb4PI0IQ/uud3E4+XNz1KBw0So4rA
eUVWuyhtYtVHdOKjgGWQoPQsN7Z7ILuhcWGM3o2Z7wT/R/kCzUuq9pDSkLZIHh2kZ60maU3HQiqw
hm3nQk6eu8ILhKK35jHOtSfKa5JgCsqYUxYPA7Dt14K8xZAxIcZsbb8Q8o5JVBPoEdnf5D6QHmkV
onEsPLXWDMSME/7nUVpUthQ+4584AW6YtQMETE7oNoDHfQ0mX71UDkYhTiMU+XODKC4h0nyOAIrz
iXUfCcWEOUURUBV9Pfzpr2X/eoiD+zgifgYG0Wd7VOUEh0NSH+2SjQ94POS2oy4sUdBH3IImkjQO
H0dZzS1LJUToGkr1yAoop0MtDAAf/KN0897sCHKM6kHCx0hWY7JqMIUCosU/Xx1aZcWGD/CmpP4+
HweQxINNKrbzhTmbbH+MwP3KO23lV+e454++6r/oeoKJLerDsgHfEZI2Y4uCVJMGwNxNgd4Qwl81
izbfKAMarBNSeLndzqLrLOwuJ3/oX/XptVwvPsR9BTSYE217creYH4f21yu8cSLzVtoMhYeTkLXx
PgWEQCDNzTgf+hzlmEmT/0jUB3Oujq8DlvX6bwlNiACsfDxhVXfPL8eAm0YcLht+vqWKMwCxVigv
UGaJ2hvbk5VK2dBznvXb+oMeDUOIRKU8tYf3gGo4GlIfsiESFQaGJQIE8D16aHG8FSBX8FDPN/XJ
KssqppLPT6qhlte0JqAvw9QLQJJMgpOxlw5+HZm0Mib6ocxXeLFBzVrHXkoZYJntU5DB5rDnBCbO
h9ZjiVTxYeE7s0F2X+nqkQYmz9Abkk8fu6XPABM9kKBjrthiZjBlrnw2OgucXSbA27Rr2sRvkFZ9
9QQx4KdKaybKlGsbYgW6tIJ/GvvhUNzhiOKUbc/19p8oNOeruGl4JKGIOrXxVamiGlBaj5dWdN7F
tYk2OpxJHSnJkblLDAjdVyCOl7QErRl3okKWTmstj8Vhw6rjJaIxe4/k39zOnC2ukVLLdoib0nWi
pdjLAamVJUB31eraWY3+lkb1lZ6Dv9fBcLaGKg89cHaJRAsquuKiqwD5Z7eYkf/7qWrGbFvmsg51
Wtf/aQOhyKyPueEDnrFPYfmiDNPKv+eJ0QWYAfeOMihr9mdjRhueWl3vVZcMcgTQfkYoo+6DRM3j
fSNZHwVCrMo1nvencqQ7eAgFPwc9e1B3oVvpzElqqI8UR6wiXi0gP1Sb8xFIVEo54QtVvgWEqXZI
9nqwUeoXbv66xj1xOGR1OGzSx3KaNPHeb/l5GuGCZ8tgWP0h/GVZIPxJucu9ds12FM0gw7c0tJPT
nzmjYunkd9ySrGyVkiyCxptKas0qri3y7nGN6yNan5IsX+duq0fmjxaPBvJGh5OEEmmlIV2TT4xh
7dhBD81TSbxnXKwuP482HWhy6778pMDSx76YSHt7EvyhmqnqsHcTr7HfeGYgUqXAsWPmq6JmfBdb
61wPKhn/FIsM67QdI8E4DkPS5CRL6Y7UP0qJ6rxl0KO5KftnevmFzfXkijMnesJCC9rhf0RNpK73
c5Z/EGo7o6a/2u4hQscO1N9wZhYs/0Iaw7CFhbJZW5eYRGGAc0jH9l3FNNW2jBa02IsCsvhFGBj8
GAjgsYPixrtfS2Y8xRfJ9djK3UlXDaeEJHZQJW3cx/2F/CuY/X/2d0mjpGA3oeLiXszSWPFSCEzx
d/Hw6bXXMf0uVevHBc2wNiSHWLB4zmtfrazXLp3XYsZeXtfWiW37//w0tjPOSPfLMCdnsbHlcUt3
YWvuVzvksXr1vLMlgzWkLoShYNrixXyHuqEWFan/IGJx+4e8JyzwqVRsldYDzeAd7twr3Qx9zjlE
7TvuhrDPupYnLBZTpnZ/FQYIN5Nkb8aemfdllSu8uVAMK2zuqv0hel4j6wpJF2kf2ACNhDK/N9q1
BYaaa5vipguLHLlsUPiPjRNdV7kHj0stkZmYQbmeLrLwN0UeGutWhnu8rTBja+84CskziePKRiUO
QQRrSzJs7FKPERobFVGo4z2wE8b28GrwpLKpHS9FOzwpDdZ2q0ndXggsA5b3N1Mpm13Jh34QFEY6
CLC/kXqtbwrtLxAtY7odb4FEKvmqa31IfTcO4IfkcZrc37vSkdoZuXdn1OfXXDmKRV19Ax/Em/kU
6f+jUIiKQ2NjV1kiI/tVL1mWFiHooXnoYdKhpMk43+mS7GKSFcVTxFKrV9+6eQph8qEuMOmsagxM
alRV3i/OiHZ22bCstm7NWJoXOJB4yDm4qSJDWuplt/YulIzfbF5QTnXePOUBbWhv405d3/PcCOo5
07xtWzlS07a+3wQLQ6j2JyKdjCbQtLrKjeDeTcj4M2qF2/22/BOy07gnh/My/kRRhx9F+73/WvxD
6KlcunjhWx9xs61lDXpvEZw7ZNq2ieEilHZqf2HuRPBTeluRCeYmNv57fvIND4G8Xag4kbcN5d0W
0JdESQP+gm/dV+iD3IirT/0Ljqnc4j/VEs2Z5tApDHDTPS/6vfUgILT2r90+EOUHJ+svUVc0/SDI
TQsJ6+QzYdFfj4OUjNmfJ0qjWNo6KWsJmTRGzhaSnLzTLSxlTojYMIzkbWIaEJQL7dS2qmz2h7e4
pCZ+tB59/wGkr+inuBBn/F53O5YB5kfiyEzDRXP4R5nCmBU6D5uaJ8FYJbY2d2Q9SsPs/hBSdIOM
h9BFt9a8gGLUOeKedT0hkPC8s+EOVc5/4KDqJBTSm994zQvqpqDFtasac4Se5m9nhyDBd3UZ4WEJ
vwG0/KbhZjfgwo0KwyAAy6E0thy0vZyZY9h0hKZvmz23Ui0faVdF8C9yO6ZCFSUkFmz9ObSjg6Xk
Qqhc7hllXOGuzFIHt2BJGVkv6Gz03WSXLSaQzK7M3aDOCu7loN1odinRN7oglMhAf2b+tye1kUFg
pIuP6q+F9ExFlDDPdNCcH5nuOBavANhjebIy6QL7jbz/3wYaVvEn8aX6JheglYnuncHi2HmWilCM
9Eav0iNE4/SZzuF0HAvgHaq4azfwTIb6/YaB10Q9VhiwhFDDHJeadfevJTl1iQPzMsDBYV8KLsW1
o4IEbEUywm68L3z5wfH0IjNgmc8AHuSgr/t3/EKWoHmeuPR8yjHmC7dqK/Er8+PQCQhUyJ05Lq8X
L7dBRXalCcPI8kA2tAUEeXb4SXA4IBmBHrIoQEH5J2Akc9I76yMthga0FI/8tiYDUJqC+2lOf+20
6yfOCWjOSWt6JKb6FZoRnbIkdkMa2CvfvCGuReIvtvzazGSOZYzV0SI72yDHVzT5qrfM4YTx0wgl
MwhawqKIqX+rzAyi9vviKsFCStaKju7LLXR0mnC+MlFkbMLwOAFZt9UciZz5ytEhWO9h+OH+6EvQ
QY2X85yRGJJGgs5DeOmtqTSqwLi+EHBka2lL3Bl68dbAwhbPQ3TH93eCDniuNitZdeAoFmoN7mN8
JhdZ+QC0C+TIUCx8x/wRVA3xSdbbGtISCzxRDa7LRgDMXVurOxWiIjBbSWWFiP5KStgrWPE9eFCy
CcWXSDIJPis2n0EfT5NXgdsYrQqsjwNbNVQzKWfgipaUraZuSPU9KAAPtk6MgPOTXkOH+azQFT55
VbvPYyOpkWaKe0tr3RsOuAgP/y8+cYAYD1tJfWl8aNXnpW5OA4GcnJvWI0Tg1qZhIg6Q0zG0SeNE
qUKGr9MQB8/S0RqoL+YIV2aIv495Zk+S7iJIz8UbHIul5nK6GQXGAMdkats2ANCfgtdKulUdhS/O
AGzCUKhgPCwSSpbhu7AcdGMCdJDTDRWgx46DkPlsR1dygCW3WkR0k0afjH2DWnjbI0k5d3HIGmK1
sO7VAAw55SNLzWvkRAs6HcLY/1swtXdkPll1gjDXENHxLAJvTPg6AEcKdrvvvHaF7xqwcelfYa/Q
jV9COnZdo2d/ZbZJQJgY2xiHrGnLll2qYutry6/XLZU+QHmj5ixHr3MH6Pt7DlHiRnFOoz1qYGRH
BiYN7MgEA9sU1JuTkiw3WgrtnOBd3pEW1VyBmwIGK3Q/bu7naTXmdL+u3hIygVn8fptlFatptEc1
P/lsO9RbwtUhBWyDz/e4TZrznr07N4KqgH2t+/CMdbTvNZMumxMgkGQqZIWQR5rX2Rvdd8qcKy7u
eVty1wwxCCO3VlN3wQrcLqZnt+1/1/wZI3KdfcnYDDtjLuCAGDwJ+35CuJ5ioQovuLuNFGQ3doCP
EyRowysaX8xZlhMnYyG21LU1lMg6nLNAFaurPyQX0py0KCCt0JZshR6KEx8hKUKqkqR/aVQOSQxu
L4qG68eY0aptOnzcziJa50NiMlayVszE13QtN2OA2rMBN7N/G8i+BwKAIEf217Et2MLudhe1P3Mf
e4Q6ZYiREzrCznfE/idhzAtHlfEiH5OevrvhGJ5fW2TG5JJbAGmTJHXe7ouZNq4fZ8EiWCrD37Ju
BVjIMt6aiG6b9gbhFYqoHUQf3HLjCPbi1VXoMAhOrlAZCqB6M6AJZpbSr2gcg2AVDDKOyZyFStHU
CBXIaTWCI0Dh8z40nm6HUPqXWRVt9bVOtVtjOeqkBiw5WCWuW7GToPqcWqGK4qSnByIV8SK9PZPc
g5jy57V/srgGYvWt4/85W8fYHjlzI59RW3/63jvsej+KI03xrjEwAvfWaCAsHpwOOjwGRGKFT2da
vZumP2c0YcceYOfejLqxGYZABcahIa3eKwudcN5tpnc/eX7ZqLmtQlKQjRl6esP1fwIRx1BYvJb+
zZJ3q0jus5SUJyUPPCqbC1BGtEO8PDzngRQkKiFLMCA+NXuxpBWEoTCapu/xGE5oUD0FgNmS+lGA
gsn3PWYq1mfBZmyx+eRvy8Mn+97y94Rddu8Gymar0gbYQL6H1h30G4L0NYP1pV/OKpTy7LCIDPue
jT1MksKN/ci5yCETf3CyQhvHBHBuFel8EbymQkNFVvZQL8mKVDjjHClt5PHtPsyCcIap+nh6XJdx
za66PcFXkot1+6MsHOJBgs1hDoibOb+zetI+sJWa+XAWVOMYz2AV+dfWyoc00o6ZRpQWCtCqpHZM
C7Hb4owYkqRSL6eksmecWHMsNgAF8JqTPsjqsyLUbPDW8IO6t/njHypI7t7ZjEC1UUh9XuZtRzT7
03rciIQE4E+GfNcGpYNcnHVusgpKC/bJONnrrXNfhl1vnJU3aV5kDbN2pNJtE/GZgcBpTw3yQFSt
22CU6s6vmsqqjjUHcoJ6UvGnN8D3qlaLS5VeU1Ar8tNXvz7QwjCQUFPDwvJLWc23lZs0jIwPLZdC
FU/gVWidwnr7fxFCz8m6Z3XentG3lJ6BoPamOV//5ZDWaIlICC5sSt3gCkKvdOJJdFkZOFOFH7Oy
jtLduUyrGMxWWCI6sLRDgklUKUAPhumv8Yam0aa8QHTE7Y2tFqkrjmxo6uNmx6FCpPKSRcaG6JLd
s+CdfgJWD3ngdwtSB7NFNB24E7VyWdnuA5835Ko3mwsQO+3nmhfi2oEAWs8xJ58uTkY8xjpr2mZX
I3Y719RMOK3Jr02bKl3DDpiRq70pimV8DtkBaOO3AJBfCQ934za9tONGGxopfrcbo0ZSzgpgyjk0
a3/O+fV0ADiiF8m96bI+aX48QcM8dfAz4Q/Ut8v0WIAAOEQdhi23e2NPKTqs0z0noReiTvhpeeDw
oIlZ3CUuv/8BKtSx5+4GGybBKZIEeS6/TWCqpENzC3RGm97zBxbwDPYjNM/ivdjWrrQdE14Wx2K+
2muMWyj4oii3mF1owDrs2UIL4+6WoBxT4dEALTpQYAdJkjzGEwn2SDw3UjHMztY/rzx1OJ7PQ8yX
u5UYkWXo5DN4IOwj0NJLfPNWU58MIkVoVDx/6GJNvX25v5s+N5QJU8AUVkNTxljPZR+jWClObh+v
xArbWRNdFwt7Y+4IQyeWcwzk8VCOjReDbJqgPlk3axdRIAIBuAZCxTe/5CYVaiugaxJxjHc+j4ev
BcsrICWebcUFNExYAIDYfXsI7nqVJAjRBF9b4Wk4tJZQeDkExH4kkL1SFMP/N791bUS6DHJSz3AG
yw6aLUSev0KiJL8K4s8jMDtDSsULJSYAgYubEkRJl5cnAnoO/3Oao7XEPyGAmSPosP6kwReMm4Mx
3tGoa3qQHUR6RMaLG9MWEJ47cDm7e30hA4i5BqPymAyh+cRqv7QNV+bqwlLN73Y6PW19KYZvvVDh
CnqD58lSoAy0yYfxfYiiSI0+Ah8gojDTrpPrTDDPM73mCyu1jixm/nlbZDH9hWvbp1rWAeOozeST
sp5rKVk7DXQBzS0fPx2jA7EzKmq5jxWyA2BVcnjLi4Pm10r4FQbgLh0v0rjx6RM5KrjL97HMGX5E
3+L2y0swn42bTBCc0NtK0W1et2PpDADHbllFfcjhbw+gyvxgOUW1EK8zLKF1Ip2NBDJ1d4p9dBLl
J5IYHBUdWS0sWyxRxUAHQh70Ya4oayTDBS5SSOCdz35UyvXb0gywTo0G9VH3QJCZlx7To1dcA/08
z1pOAtLtCBBOBMj1VZwnCJoXNmRWT+i2MRe5SpCiZKvwYCtVy0xpw05d3/GhezHpfVsAPvHAisbq
S68cvg8kRjq23+i2mcDiiJAReIgyVcQdxvi17b0yzOTIGerHN1/yhRySh5XZdEMHjpiDwXIIfVtP
Fy0zqrEsFdIQ10GlOZs1WoSHh8+G72cuGDiGRk5xtwUvQkhUDNCYLBtty4ubgzNu13arTXAOmdUT
h6esTMzk5jjZMARiW+kIMwMtoKhjHPQ+tDAVe/HepzsncFOw8aen7vbGfjIc4ZMqTK+lgZpalSoV
6MfwMrHDOY++BaUDCOmPZx1FC7KUoIK6BV55K/KdEW+TdiLYcNal9si9CDcaoMcy36wG/05nOdZR
zj1tWlqg1DJz7yTKshY66TP4lZXKzapd7xLDfMjGF6dmLOGJKPGE+TwKw+xN+LGZb5W1Tz9j6e15
2/KV13QLl/1SeyHLGHFv7ctyJI9eKcuse2e74jINxP3nDSylNClJwhJxVC20lkOzOvM0rL2oDf+r
BShn7g06MfQiYQAIwPpazDD0uk1ke5IcfpsRELeQEEnXow4ImQgmTzqjQsES1kBx3G3Rz2VxQ4GZ
JSSZT2HfL+Gjiw47P5HP6d/VK+qrlATmJso2uOech5w2k7+ucGj0kfEhRh7rqMVlHz54tNXNuGTg
G4j8mY0q/VyTXvXEYyr0hhnrIx6E4G7vWvFFMgriHMAQ6MWNB+iWkFlWXKOlNbek1BsIw9aN+XDj
x/lqqA2lcTEn13qzxKEzvrzhb9rc4nhU8HdwHq1SUELVcrrihNM1fdAiXEWQ5fgJSJFxwK5bhA1T
iR2R9cvzF0Lom1EIkRwQs6SzPsbdxe6mltUmBcoauYUiKiJqGvw22jNzThFHYMRiowDqLhLgZmS6
q2561WdYKrvST4156lA4/y5MxHY6dnHAu0SXMGcCcYeZ2V3zeOGtTb5m6B1gBRN7bAee5DZOsjg4
i66D4K+/O7WfeX9dD/fKFMqmwVzJp9Uf9doP/caGmNCldRLb3DnQ7EVtNC3YHUD1ZJmJ/xDKMYfN
HdjP8sWHMQHY9rKofwg1MmssvOZekbqDd9BVqNho8lKarGcMeTfDksfxCRUlYhhYE8r15uRIf1H5
CVbV3mJmIszksFeU7jmZJ/zRPLT4K1C0kKVEXb6s+cbSVyzgWGKftENnKgTDg6QjRiPisuZ2kqel
V7U2wQZc3USbRZUflVqtbuimZqClPGNXRr/haMqLwaQAy949hrU+0yTZKeCgw8p63jgVnwjD1VPw
4oxkzukuWOIx3J5nxPPTH4uVJf2fqLUo+INUNGgkaoWDV4EFC2rB+VRjxj7ng3wYCwJKY+mnE8U2
ds/pkjsdm02xQiOl06ZutMlyXPBWVremqXObZCM/c0e3wyAI88M5gL9qTHEV3Qbr1HMRaiJprIxb
qhddDRqMo23LNv0OLv2j+6p/ky2n/A/51H4aOs95eZ46xdI5A6ZEcyEVEld0rTD7QveNGONdD4U0
xqs2eavIdbSmNgZLm4hnQtlJPdk+u+52XCdw8U7QpQ1gn98f6HMrywFSixjnqIaJ1jp1hfdIOtCx
cnJcCfztjgjlkekiyx0skue5hKjgtpkhkkgMYgGm6wK4K2bIiLTOvJ7VlPtA4AMy2EmyK4zaaxqp
uLY0ApcDJIQkGvsZPxOX5srcClhGJZ7bM8IggPkY22pT7iV6HHoCKHpztIWaA3fGiY6msAq3dfyr
H4/DzvMJQv0RttVIJSf83WjOd+0rioDhoL6jWWjIpZTSL8UwmbWv/HFFZALak2kNKY4vPk80hDGP
qILWUWGRXSCrQOGfvRra+nRvXT4fjt2EQ+c+OTd7DximRSoZTMJ4JcfkMAi8/JE8qEZfZl4QMQs0
6EQz1fkMMVTvbwiPtR/fY85LCvoIzZG/edY0SoCU/1Iq/QoTY/pLQ2hpHopoWWQW7SZjqtcM60lN
h3wW+sJaPE6x8Iq0GWd2qR3GmUbyirGK4YJciJjj9H1VMc85ra1deiTQZl1wdJ9SoaPkcqSFhCSh
aV4vCalHh3d/g9iKEhLVgpfAbb9zpoe0NeSJT5m2pAP9UtIDpvPmEUdcptwZIY1rHEX6aOavrqgn
eXuv88d2/cALEwnIB4xMVff7XAgTyEz1K1oE1+LvXKJ+wg1Wt25VtR3OLHLDFj2jCGPxkC+DAFPm
qODcs6ft6BB8+G86rzIWIuOLU/5VOSTOID+8SX7wipEyXAbVgzjYb8lJ3VdBf8AamchiJWcJqxVF
/88Z8px3oBEOQAuM8zQukhAUFDsIRCuPxrazKpiY8OuarkaMrGdPD3LrItEmrrMsBs1YH8q3+VDV
w3zqTk7aH5cek4jh4nQsi2eoJuDD95B1TRy4y9IbTzxPguMWcEpTQqZvmbZ+MWXWmDvfDApehSua
Zn5Sx5UBZgoWXZhf4DQNWifQEMWmbxxcmAf5C2f0xiGbpbQwtiNJG9dJrzDbcU2/dTXZr8Uguoa7
30BC7JJ/IhNx/OaU+T8OyLSt9f1iPQ8hreBpzs68dkZjCZH8QMKhDdtfyJ4P0wMhlB5FcpPcqPag
4wcsm0ec+PmauZbU6nfeN+Zc+ox8K13qCYAMabuI3nAj/BjIwtoOY+Os+Re6d5xwui2gW4U04/rs
Aex8IGifFVh8ZBBpPsl1TKEnfn+gtT3A70b/J2CKu794LhrK5EOr2yGfpvjLPqiCfWOH5IztBI+O
7yoBHR2FLelHWc9lu1JzH6JQK5ExnhUtU56MW329C2uRqOMDZQXcZugS7X3SpdyX4dhcZK0FgP9n
VSpK3pWbLZ9jGUBEYRE7cPY0jagYqN3yReenIJLZAO0CSw8zT8a1jZSxy6lwxaPlVFKbCjedAhC2
e0NL6cMMSEN4b/XSJRMwrEuBZMTAgE5nx4cGN1EbRUOvwUEVv8tRPd3wq79wHdGWW0srVe8Gif9+
PAaeENurunH5cJdpx5LYwfI6s0Srrfnx02YdLoPERX/W6QS65BNp11FP8EHQsaetuAsXf638rzKK
bA7hbMXXPSNCrBllpqxpbPuywIghxmuO2dcdtvqqGti5BbADxaA+W66EIDiG5ZGJ7nts92ZWlgL2
rMT8/Du29ZxxWjgGe+VsYi04pfKgFS6l8YYm2AAfGlxeQKUeIz71tt7VPLLgNessziFVyhFyrjl4
9rbi4MyorA0KxC5774SKuvJ5BRDzUTV0LoNWCfV1AgMAHDetezl+jTb96L+b9YiSdD4R/AEQtCQe
94CsKhoJS/LPNpl5p5rcBAGndyttiV+9ytbWTHorEDLAauSDP93Hk/JDlqcOB2fxgXGchrPztAeR
V4ypNWTzqrLp95jRpwH6PQryfvBXlk1V7/Pi0HOxnXFe80mccD+bUKAMCzZXlpFrpBAXEhUG2ePO
LaDWgZ4aZ27WXLUPon8QsQwSKN+pUIOK1iQPncxjxNjOzUAG4hI0ZnLnwsAdDfFqdkcO6xd5bEW2
+QQ3Xz55iVef8ntE11Csv6nTX17FWfyCgSvQl29XJdIQhnjN0uE7txZmrLsMTd0ME5dv7J3p+8Be
Yuw/3zbqbr0gP9v4eTRqyLEUoXClieIWA+S7f6ol29ktSeJz1jisrozroV8=
`pragma protect end_protected
