// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IYpRrT0veRZovmwctbCdz48Ub32dF7qRpxGAC7R80580LDxBYbHuYLRfeMIONbYhI0lTxytflmIP
yebSqtTjR49m8W5oDhLg+uwdh0HOdkHnNB54qsjcKFB0YlpQLiE6h2F8rk2JNiSzDf6l8bU25mhN
9jitT3JSUap8xiDOG1I8xjK2Yvgg2B2QnJ+V0UYYhzpFnbkVZDEOKsExPtjqu5em1up7vtYB4FZe
mpg59t3tP4OxF2FSYkaxEKlyF5H2t+ZkKZu2DFV9H8MTZjGtL1cU1d+MOUN5TknomFR5NJ7hhf8J
KwdhDN4K+0rakCWahUrHkN58kxJ9qz5Oo7kvAQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11072)
n4XO6MdJ3whzePFm49TAFiZbfNYoTt8VWax/f7E3fE72r8gYBeI1lLpelNmqlAy7BA+dx0jQK3PD
TLxQAtm467EzDY+XnPfGsk8ekQobS8++O4jejZewFOFFrDQnuxKpSvTiMhvGkBK4xjvjQtV8v2rr
hfwELBGBujw2g34A/c2oDwAP67TyzfiAy1xsREuqE0myn1rsybnZKBuC38uvyIWnoNuf1j6AwZUO
E3oWHUYzJNXyKHyg59Yutfc5ej5Qd7Jw7dGLzZfQuzJ5BjwoLaokFX8p5DN+nCauDfuZ/mxGMoi+
6S7atXt62DvNLYR+w03JL9nhX4CKpgjawxDPVdZKofv1aGk1AKLoMKF/DiRw6wslzXnxb5tsYRlF
gnf0+HuTyTOf+zcDhiTJGMtoJojO0XPuQeRt+RzRjmioUZOVQOENWFox/XTO2MVfkbHXRO1ndgyO
eLsjEFEm4+AgZAz8KvMLdr+B7oNCWp5bMHgrf5BZqU6EHwVHOPRCVDl2Ha7m053LbGZx4wiYljJo
cTl/TJDrQco7lO9FNKWR0N9z0KZv+U0RSt/060Ep0tzdBHxDA8eY/s78Al+GjKb5VsQCy1WaMUF3
spIyq44T1WSWNr7lJdnWUJS+/lAfyukB0xScktcdjdEzfEDjLSmYcm2iIKWrTu4Cfo0wsKG0EgrX
lINAL1y5jNc65yvDhi+77xcs6MZy8A7QB8qbxIZxlevRuaZWLzLodUJodHN9Of+1uIHj68cxSvt/
a/2OmmC/4umlTxNrRv/lklENyDSsiy5z2FuI86AM9lJZlfCKzZ07xDK9dpHO6MsAy3RvteHAuoHA
6GpJovfCcjF5UmXm+x+4C8w19h5J+02O2sxBBtb9E9/9EJJu+AZeYDWY/Oj9Dbl4JEZre+YvMK/X
EJnhoFRPT1/UeKjCRYtr9YyA14Ubkugr9U19y+N3fezV+lMlY7ER/qu/6gng4JUv/ccScHrc5IAW
iKlYyfdupk9GqlA/rHI8wCGtchK9mj3Sa0wV4MKGkEC5LiwxQAYZB7rR62Fedb23ea+C6T3gS+zM
tKnAAEIdq4QsQAmixhkiAYFnLdcaYporLeXLUEOix2FfD0ZD7MF3awTHhAJbp3d8WXCQAS5bGxhS
qJ1FO4oS4M39jrmA8g/yRIQi5RKMI2tTAwcGfoX224h05iA0hlHFASQjxXQaHYzeN/hBxjN5SbSj
hnSePlqslk1SjeBSl9qMKS2lX7Trh4j1wpAsvrgT33HLxHk/HKpJtUt74UIjjrF7WUqogrBtpl8A
g/2jy5VlAbGvMuVHkSoznD4dTqHwk/PjGUY4TlSuU9j5I4xj2IoxmkVEbbPuUbF7mZW/APfd8nnv
6xj3ZTVWjG0Hc2Ypj5V0Iv6HHTHJK2rWSMbU6S8JNJy+tNTmHQ4UkfSvHfw2TVpUWLWORDFKDgYs
/W2+SU6U+6CEJoDw0NTQi+iorFtfNBkK4G52oE22/+OqU4PoC2UEG0HGJNCuEUp47bly5DPPCGzz
7in65yF0XB316uk0v1EXq1IwaHtvLDXKI+l+0D8Ul/JpzP1Bd+Qfs+8ZRKiWLpcwIQZ5NvIcEagi
8ii5t5lwNPgtasR49K1KR9WleSlxJgiNR8ysLXxp1WcbaUis35H+YY8IqWnYuunD81tFRWePJdDB
O7uCr76sm6Wvqvz5tnMvAQ5M7YyadXTUw14nW/M79ErC+Qqz+xxtsDwcHQ5PsykfBztJhu5l2pH9
G9wF9GxmZFmIbFDc0iZEBCizpMhd1DEF4Pezh2rd99U0GdSCfpcA7hJRrvM6fh2h+06P64HsQMG9
zAbzTg1ZGFBsz1Qzu1DiVawEX3SYaNxo+sxVEv4mFXaNRObyqLjIX6WVvdV4qUHbB3IqAFhXvu4j
TtK7cTQceN292717ZRok6ewrDFTflWWvgT7rQeysjWjSKaQEsvXUs+BG/+/hOEsMbqlQka9zsXS/
ZSoxRoMYT7zHCMnzsYEfvqHjxXH24OeC+OIIxLQvJrsVVS4M5KikWtCVoLOnyJODL4OsGg1/NL89
CRbquPBYeDjYDMEncvloF3qyQG5veoBD4iG8NQWi0xzK58ngM9oUrLNem+TW9sVcku3OEi1mohDu
tq6Bdf8KAPfYSLkATXEnQBwPRnBQnTVYbY3Conabg4l9Ajy7gjNfNydjWAlREVDx8/m4N/x7Gtev
EYHOR4Iiqj6WjCRhvTsiOaimS2VKDxjZZyzBYPvkzofQv3QDXVpn55G44XmdFa2Pmfe2ni36hsIS
cb4DtzjDFsziRukLe12hwyTofRP+9dYgZUPThsD6CMVANJXwoW/8zy886j/a0Z7wgguPCYeOil5U
WFkzYS1prug9QHBIFnzLhRqTnZEvKk/9LAPSiRRC5itY6qH/CN0BDuHxC0WjtdvUOL6Qnm00+BnE
bHRLL++WBJv6aYUl3vmocX1FQoY5VfqGiDXZ9EARmP1l0qaF1gU0y1Qt+CSeU6j0FdMHEDJQchEC
cxNnc1vTVZArfrHioNBFgmW2ltKD9tutuwNki8LJtCSh5oxFU9uKrdWswnroAdoULbaJzDq21z/s
q+ve0Q6RoJX6VzDSOAo+MJdnwwsny4HAdIvQXsMIkvJ+oJbB8RVvVEqSxQrDJWE8h8gNBxOYH9fZ
QS4wwV0tR1NOXRUmZawSfs9c3KLDe/oUBhmXuuS1Lx9QNm0cMNahlRbrRFwv5fcSfFJKuZBoy6bP
1hsaQ4cjsWAOsbBoO3Ui6o4fSplseemt1ifWw6duHZtFbRafhKxXyyJn+T/CcfHRhf4hCrm02FGM
2FW5K0rCcsegiu0fL6THWi7AWAQ97xbsGpcyTQZC6xD9ZxUrQg1ol31+ZyfrtzwGQCdASpTBHedA
Kc86K6lYuRhNhFxhA9K/mObIDPQYLXBZPXoFIsE7vwtSILevY5YJz8I/JjfRLA2eIyhivEvcTokM
RpWF+SfhSprrkh+pzuwMDdqqbK5aFrWSzzeRjmHjwAp2+YhBxhPuOLbrXGv5S6fwwjujQFm2IUTt
Pl6W6sC8AYdQ+bzWnNXNgUfaXosJU1y3YORlgqiDhEE/X3O46bG3qJ36rmO7+eLqAigAjGv1bVC5
eeRTxOYS+fV0rVi7gROTkuNDN6bC0SlwNLV55YRHPH1H0OhY5mcdWErk7SmQrpYxE3QqGxt+VUFt
MLG2wCuYRYls2qjj0rqQ6k0oCjpngb1HInG74pEVu5wMjcZNPqk/g54qqAthLxVqzrAEEZdnypq6
KYVe92OYN0ACLi/dmvHeKig2KqE1pcbD9bJrUITsetTYjd5kBEtm/ToYbucUD4ZU+tpVIjhGoKZb
lVrNagdU2GXaAsXOOqxGXM3xlG3+xx354sd2dgllVvEwJqMsaCch6xrvI0oCZFa1N1fiT8k0PRxc
Tl3ndmudIKxICgZe4RiuvtCa4/YmrzC+p4ndxbrlciistKvmoH3cDxsVggX+0fMHMyBueEC4HmHZ
izKG0KzxJqFFwSO1nHI2X6O8wS0wr9PWtYBd1Ss1G+3LRMiVjibza+rmzM/hAPZYnVBV+MPQciGC
dF9kJ5aQeeBrkQ2lHLno1ujAVgG6iqvDEb1fTQZ4G95hSaYtt8ViTCAWShytQKQuDqLMh/ECwibW
SLImx9C5vSPneFwIdpOtIkMRAY2k/J1NttoS3vT+ZtZZ4jxJ0llF8y1xmIkk72EXa2m4OB/B+CRz
62tPLin4jMhkBP1TlR47j9/jLuEYElmy8+gBlGeEc3JZLIU1LCVOPNgtZ0PgFzevg0SO1PqQ3rzm
Qmo3iEwiIeL+Ij3kaEsHewtylEjnBXnyX0fD6tykLUKZzKdNg7P+0g6km8vyE1v5DoSpsj0ebsaf
P3TiLd7VonJlAK5dMpWrvytGpA/Ev7F2GELDn9xXXROT4dNmsXQfobZyXXe2m8pscqh5YIuGvqy2
suGnBIPM5y4jvfiSo/Jlh6wM8pM0HUxmWQZnF3kq0Vt+YcdZHBQgN8NAp+Rj00X3lh4XPdk9aXNY
YixFsF3PrOsvwvCeGZHRqxvl6mjRlpogTJ2i3K2G9HruocbyDFeEo/oNN7b3brG9Cqcb6kIoW+yV
xuLhdTfiBCax4FgzL39XqMCLpVv4JUVYP1G2rB4QpLPYIEVNMjPvrZCcUY/IhD8GM6kMAn0Q8tob
Fs1kiNw67HSopI9aOpspqpsLqbZrnJ4WSJMOB+4Qgk1R4tTqpxTQl7Rz60yrY2FG7IvMneUnr1hr
lx4z93tuZ6AYO4zGb01XoweJMaL9f6rhNF6Y5q0R4LzD+cRu8QiIOM4/JUnH7jG5bfa26TAD+GGx
jEM+h2mYsNZFiahALef6uayBcvHH5yBAe2o7RY7V29AQ4pwZK1RAIVbCAVfLgQiNcIAZTSp/9Rfc
fQKVt27jBApeS10RKlvCYXAZjb6p4wuWZXq+3k09kjf4hzlwxpQuTRx2x3VhXmzT3uzLjkEDfqLN
gAGgSR4Wc3poi2eZvDwiJhTpHOmxzJw8qSBWio1LssB8xcB0J3G6AvREaJXM4mcXcWSm9uwZl4Ou
TrseomYtF0ro2KydKCV+R/5gCv42K30WTyNg3R5uya/gn1dNryc/EHg1lZ89uKOnb+am++GrPbLE
fqYHgxQldJ8HhMLopt0UJW5M9DF3n9jvEKpi4UZ7R3pAePcnWIAHUbKRy1oaTjgbuF+X8kZdteyJ
TXEPNANDWwbs6iFeLjksgj6MbcfjWRoCdFnbKIWHhSJUUExa9UY1gp6U8S2a73Mz/CAmOd60AmPf
AyZqNFKjnaZ6b4L3QV3fMwKj+grlKxgxng7m6l/HdWB5YYKAbI5lcPEdmdUlU3lQ+dTO1X+rrJm/
hiYN3g92/2ekqsPZkeUCwT6BcM7rVWL31sUsTMD5dDQrORNYOVRueFL19jjsZSRYoYt/PsPz65eZ
q1X1jjVkJaDfkuJXioMH8vPYh0llyhdILNWYpmwp/H4evK2VuCvEL47A7f4R3DsslsxLUmCvBPkD
jnfvoCnEfphcrp5EOzD13L4B7Va1SAWkdIy396gRGd/0rahdm8cUTa5TPju6NEDoRl9eslGQDgnL
MmKkYZCGsNQgll1FXkV9G7RI7qbAE75Ejt6fhAwwxWjt82XpnQAXyw0I8SALRZkjP5UEe8lzHOuh
EVa+2B90YaKXnXiPbbMVXlihXY9ykvzV0PCVPbKhTSKH9s+xNlRW+YZh4F4MlbtPTbViY2OvtuZ1
7mTFK8iABc8hXxSEKR1J0wTbFQvOrxPlIDSux6vs7b/O0I0gGNPivlcfqzN9LqYgmk2lZQiQy4+M
ql2eRmKHC5mdiQhG1FxSHjMI3F2ZV9jr2MGv2cH7x6dyRyFnn8MJrr65LjuEF9LwfdjXqwCJGKfA
rRgyH8dlPIERSXYeEPNu++s4ClYtAb1mlLJqvdraV0uJOc5oZIJwZsis1/GhGJjL5xFmAKzjVZpV
hBApphYmXEocyIk7oO7kYIqf+BsKk9MjN5DJtKsdvlz+KVh9bHfa1k67Z+GaFrLdbC1seQZ7mC8N
0jVodppjlmaAYgwYFqslmKNTTvcfsKDsyUWxxeJnA3Svdf6JtB41h/tI/F8ejpEgpt92ZMp2Qm2O
gJIlltW6afbBYc+fYgBN9A3k1iMpgTJYKYUZLVPPCbD9SosEbGDIGvnAhkGOvsGrgc9hTOUIq6t0
/WHA849xuV5UfcR3Bmb5Z1lBRi2FA6n+uZzT3dtQWd667IVeZhzIVLkl5zU1K5aqM67HgLKLQR6S
eFDzLYOpEKJOUnxGushP+ufeGW2uPdbQI0wSMzPcGbn4p75JqydkZ9gKQ9EShJ7tH8M4pegOdDWP
UBXpUX4KjjuYcZhTZiBDVTVQitMIcn/eGyCfBLHyOb8BPbhGiUuSBEZxquPbJun/oatOtf1O6Egu
NqtD67QE3BQgJLVaYsCxghPg2ciAJYwHk8MZ1MSUqC8Z+Zqe3PNLGGME+WgDmEbcQMME4dUQOg/6
qg4DvQnOLTpVa5ZA0OfPgwIK0nDogUMrptvP4ouKQUDO98fCuelVxSpgbg2GXevGyrAWL1bodpw7
qmC/apYiD4kQ1PEL21HE7dwRZUj9jAK7CBoMHKP8nMDREWFd4Lbe3K9dZaaCBAy/G1HzOKs8Fsff
x8oxo/Qy+n0MwDEduhzptfM9dpJw30O86tNLFr6wXqp6gO1IBLhFz/sK597Wb2Og+U2g8V/vGQsT
UdJqB4YJ6E/dIt+mmIbMEh1k2Gz9RmdS/5iMzrV2vd/6S86NLf7LIoehxJaXQaP6ckT/tROAUYoh
4FoqSkQLNej5LvxKeCVMuK3ZhbXnbLmltmKY8gP/OwqjCUiPqm9RmUxTQ6WraGYRyI/4AWQHig57
QqXTQE+nloA5IZ7JZnE3zpJwvKBsjHRcedBeRafpd8Yc++1XtisxCXSnSn3bGR6wZ6yiyKn3wZO5
X8KmILFOg2t3R15YMdduWHbcZUoQRjdLPEtXor1uvx9GhRkpyJHdAz3a3Jsm2ziSVp76EmPOIwgU
TLdXItjHCqq0L3KuMvbDqV6wICd0ynMoHFqNkqXZylUPfwG5S4e6IYkiflowI3PGp3BNBzKrw1Qt
GMBFoVZYs+Wd/RM+ARD7mrmIotVQIxOUlKEDqwAScLYpaMi2xHN4QxAK8YDJPHgc7q2Z5itSJW6p
n3RI8gj8rcoh1Rr1cZJjPpO//ssf6tb/eu7JEkATOUleOR5bFGu36TWRmAAmtISbcgQuSnHNLkX/
AnEOeHFfdVqHFEVLyiEvIwp7L7CwimMFtPvzU5nfQ2nVEd0AA06ki07oPJGH8jBjjQteKTWxGVK3
xIkHkTA1TymYt/MLboDKQLtI39kIttSgyaW0RhztMTr0ihMu6ExPFansMWt1cbp2JLRyGvsTtKMi
ZU1JBH6zBIrJf6iV1GKgDR/1Rsr0693QSXOfY7zwRVUdsdkRNXeDYv7KS4bnxChXGjsahTRqQlUe
PRdnl6YqxNDtrLJHVAFtYYWDf9itk1I2nCbquxjWUvMLboIvJAJwZ0XCyWgTi/QjNAGozHF/Jh+m
LKYmbpgImKJxxo9Nh24y8owP0nY7joDC6Aq1isSLgjJFwldBCRvciFuP3miVimAZN0ifniU3idGm
5xrE9+Uj1KSjFJQRiUTU+4huLrFjC9BxfU1pECczUPe4CZRpR8v2XT/VIK9b5gfbcIR7RqNsilpD
Kx98wZ4B6SlpJdPRcSxjQyF4LorWneCEOplUrHAOVIhufQ6Laj5jEmJQszHSYKQrzarH66eemJE4
nlXPgL3I71SeFaOEwhUj5YTKibGlixEmYT55fmHST95/ihsoPUUCywTYbVrf4Ob3eWizVY86bbL0
kNwh/ZbeVlI93ODvmsy8wxoR7EsO22RbP32p8KwykL4BkBV0drsNuO9o5i+H50M6pF22cM+VIoJd
PxdyzTifUWjFmynzE+VUZYaqbQ9vZ7NZ5QfCXDB5EAgGmWU8N0sqKOEoUJUf0UZRMP5FwdjnHc5U
ODUw2l2nDkHN3VnHb0kc0nf3r5ugw5Kt96582b9KsTSptl2yuQB1jua1szmluhhwpR8+d++Db9l1
IBzE4UmlYCwZ0TizV7eGnAp3nDLD7qAsXU/+49hdjo25w55sIOOXsV1SDlbMn2UdvnNWvkqsyiBZ
iQc3+J5EyCa4FO8il8UhPimy/KwUwF2dj8N0CjYjmEL12d7HPQsVJrgMWHMa/a9b5q3WShHZWywY
558korYaW5dgriRwvxODfYiPOKPnauVNor7Oq4p4IrAguwKNyvZj+6ChQMcVs+AZzZ3aWdapWIyU
dYB5QLC0qzZnVlfdxjnjPr9J+2bL8mNSxSDt4uVHD8c6RFENLnkXvvWaGwn4DtK9xz+WL075ulGJ
0UBy7AqSYiptkFp/+BkJNRHAbv3+ttz/TxzA3KPh2agoK5xImVB1A3N/ArCQeM2yivm05Lwr5R1K
k44dgUxIYSeTGKAyM8k3JwVjXMUfMKZNQNIXtmzqUVL8zlsfdwvZygn49CmF/wPJVn7xsgHNUfPc
UJ/YK09Tvi5HlIr+0nCXiQQ7pa+36XPwtOPFNWDNq8h+xg2Bi+UOVTFazOt0E9Gi9OQxm97mxrOR
+/VNfuhscM3FKAIsEi1peiCBGuvZuW2oRDh3sSsbIlO4swQvF6lqbL1QbHA85RS0tRn/be5++lzk
/hGaDgm09j7124GABG9BU6r+gmVEPrQcPqI9x+sfUtP4jkrlDKwNIpvRKHJ9Ms9HH+2M1QptT7Fx
XbZ0F6GZpCkihqIkLMYfct16VcYoZ0tJFcmctBd4mhEYNONBC75l1IMtX7exsAz7RwwarGjLWfIf
n6PGrzE8PqhAv9npV19VcXnHeK9SIqAAxuiHEqaZ5yw85pKXekxt2hGKTEya+9BUuHluPx2Np47q
fq5XmOX8cmdXkppx5bJheZQ9sTvtQE49bI4M/RhvWCcFtWmpjU7WvqJQGtDr3w8dr8rvrDTN296L
zlKO8vMzgyPYKIs5qT3uSvjWG/z+JxMUGrfJ4F7Z50iOlZrpPd+QYC9+nZT6u/yv4155BC9Mvr+q
s84pO/ZKIlPg4mEVwDaaRLQT8AlbCMCRTacbPuhlOpNUKgQeOmfuZJel2JxYd0LL1ql+KoZfAKgC
lrUS5kRcFyIOMwR4k5oMyNvea7EP0SLz3q0mJymCX1rg84GTwmov79OzIg0lQyoMOL/kMCf6+8/J
7sX4lmC6SWQw5/Ert9B3Vpn4VcsobJXyYKIwYqQVlR5LIozOaBGIQq82KWHL8mZbjjMXvlszt2AK
+sibp8jYQdFnRM57kwz/XQIS8tVP166iSK9xaunoL8XxapUOV/ParaL4PlfsekqaBmia2QOCjLFb
PNHKJ6+QjOwcdVZOMjRjY/zQsKxaO1LAaf/Vt0p2F+u+vd0iF/gk4spBfs5FQHKywxg+f6vHKcjB
Db2XXTYH0kURXxNns9oEFVHodK29oMdtAoyPaD7y9fHT+2qwBi9bwCUK2Re22bXX8487furC/z6/
aaXL64j6rZRr1oxcFX8Al+kiaBWwsO9f2yIRyLQTOpgleOTHRY3fR7qzz2emwDPCR+7VDiV2a2tS
eS+EL5CAE7VTLygah/1xGrGqDhFmq5kmNBLztrykk+Fsrh3F9SICE9pwSpzk8g29+P6YfH08vFeC
QrGNyx1EiqZn0m4wfN8Dv7LSXfCCUGMK97fb7YjyMJomA0AytbK65oefb4JArDrI0XecVW+5HycA
syvg2YtPGO9QvmGCztWDV/hmiL7UIuLDnYOJDRVkBgQOPtL/FYYj3M3uEeN4XMc4u8Jdfa7yxkev
peKA8qzZ4Y4AtmhrkrrpRH+U3YGpknzkmb7DEVuAre9nm0RV6WPfTskpK0HjSwPL5bIPZwPeVLfC
mLYccMe6LLeEUc/xiv1eZapHXxBuqU3XaQ15thR7BisbIrDw+F6/PcL023lvcjuvUmi7JpCtrNDc
N2R9GZrwYH7Qcw7luX2awHwmgS8/Jf64UNB4nCy7KLvPc5scW5DpnYGezmLix/R11TJs7bgA71gu
vbnKxG7XkgXyT2WRZtTYSTwKivNhlqZ4Ql5Y21JQHR1Z60uEG1vFZ+Jms+lfLuMnO1R0sYaaI3PG
Owr3okA4kRd64yxrSvZnPb79eLGvBhvHr5cuNJl93iJO8PpBxm09L6qcj6jRfNgxQITLKtVEgQ5F
U5EZ0sV5RvTm291oTzuIsovAE+TVHYlEHkGY6qCA+sWT06bLskMwwz9mZFB66dLikGkV2nf2rURN
f8NA5/5+UiED3eaXGJPrnViXGkVleyE/YLQAhHw41XPZSwOSWmeotSnbyJarIPezTSC+KG9RGH+h
zm4hoK2s1j0h//iinn7+z2DHdj2Fri1A85NH/Kuxh5PZ1cs5Jm/Ir//9DEUTqiOM/NsV/1wCHHfx
P575rksIp59//xrIwQYx/mI3i/whVOF9YZwJX9lMFQNRiNt6SI71V7yeE8FGJatU0VPrzjUO/YKD
hZui4FQ7du22mAygo4mZ8+Xl1JQuFZW+SCiF+26yANgp7hL/wT3L5lqb8J3bx6b2oG6LlOJIFFjo
sjgmdzl8zbnX9PzR8wRmlSv9h06zPqe0q+vu8H7RnBn4WYNk1fJ7auAtMMH1kiXHbwG6EdyejYew
ZxBSevBJXpxRG088n+809QqqVHkdLAnaUdFNf0tBql9GhKWd8qUT8EChaBJLeWvOSk0myqSAIENd
vd5v7JjIMw54mSP19rMkHvUThzwuCJAb9GEjKX27xIL3SGY987mMgIz8OwCd59DcydUTIskZs9qc
gkiYOYSiCN8kcfC/3CQlCRH0AplNuwPjBBupxfyFK8CPlkOEL49DUmMcmeAHyCxSTLxBmCMyVIsY
ib9kIA3MuWQhk2V1kpRySvqjeb3PSlWXoQpVTPRnIGRzn9hjlC5hdYzmyZ4iyYKZutIyvErhJF7T
Gwe+WLzm477omdHv01wowK2VatGCZDQLvkiCcJXmoioLe7kvLo/6BA2M/plY6iMHdRfzkxwh53l/
7geSZN7atTKJUKUZwSU9d560PNzaKrY6DjPrroXQ6z91Y9fPOltIrYNC2/cNYURGcg4hBsmWdtBF
cJFZWUyxZpcYffOh1ZlnMM3fPaPJqP0unHIIb0G3HpU1UMwSxGZjBxoOf8II8u8vOj/6l6igp2mk
xspi4YRp62RUJcfxhqUVAUUYK+PntfQ47HwEM1jXzy38jIlPYKaKzAAIuKoOQT6utg58041mIdSA
whVayqsN59ujG3Q9QJ+DiV0XatFb6k4AA/+e9XOyKqwgdsxpTK0ZZNkYzb7bv5kpjGQhPpPcJBVe
BwlWtG8/H1WEwKzMie1dcM6qd15DBR6gGpx1GUWu4kn8x4Nz9KaAbu7WrLCa/85Xen/0R+6XRruc
kB0DSFi53FDTiGalMByxumcykcpu1gQlzzDw8I0QVrDj4hAd2c5wfUN4r658EQA9v8XZARDSAedR
PfE7TU2VyeapT9vGYdhajUXGksbN41h72CrqFvQ32gN5KgkeQAaMIoqMxdfF47soF0LsLcfH9RLM
4MYxR4RcVi09zO8RxBHr6QcTkIxUKKISUTnzG8zjuuohFCkNksgIYY355IDRx5OJk4D2gdNlTWvC
cgDc7XLvldVCukNB3BP2BpXzA2qxopfM29eQja5DDCNfQpeu9Kc7tr66PdqH++qG6k90iIJXF9wI
5k3V5ggfeuNtnY+GPb8USMdWQCY4gj2ospuoCYdPljHx6WHW+c0z0D1ecsS+MfBga/z+CTJS96Xj
e09vl2P2qd6t6mAmxT47hfaCtI1dTS5b4hi8r3bVqZao/2RoZnGIa3u9v+HDjHSnCGqx1RNJ2YQ6
b0shnCPnS8SaK5qVM7j6gmW/qvndPFfViJay4NmT3dugm8TR7GvZcIHkX1qwWCAmlsHFMgCiBacR
PfnFa81nkrFVlYS35NRRlvtq9QWWUfA7mQ7QVB//runAUzcoq8unKOzdgSH98gM+Nsd42Pqv93ys
tBQEsmO2ncMVcQspNv/kOpUuqJDS4+5OsTPDjGnKFSj82cDh2Ia+Klu1qgau9cYJS+mmCASLzB3K
pXt60CTlG8ksgi21H1lr97eJI8kksuU3Z3Ufs+H/oURFuqeOt3e1SxX2AeGfKr1+KUAqtKe9dois
C1UHr49Brbi+0NyTz2M+FKUfbbWCLTeR8ymIWJAEeJVOJGWC4DtOyRGNsaQDHNqQm0eBNyd0Pvow
KWWfZ6PYfKuu42wUb2Xadbp5FILdPRZICqDHijce/YTasRTimdtHePG7yTzXzw8YvF+y7BDIovDo
ztG0CNk6bASksjEDV7AE5RAlLH/8RFEFEC1NXgL2pMWctBttpSQMd/nc7ShB/7+ldVZEvg/5iQPf
Geotpo7d2/QsVZD8RJdobkdc13zQK9rsP85u9wShLCOVKpoHKPWg3wmgGNIhrwL9VEfXlOmjgwzz
cZL8gCNh0oNyCA3vxAM7fyn3NPj2KImKoRoN6KikDCguOYYO3No8wd5xnPGk9Ejyp8sx+k4hMUWF
u15yvhAo9IrPzBDWKSAIyImIO8PasmgJK7GTGI3HZxVU+RW6petbpwsGQSjT7o2jhBVUBhjfaHMn
VyFck6vC1Q2TJQNgS8za0KheBpehjRyI1tbsb1rpAPdJBtj3L/PDF9TRUooK9eAjLcTeyRBYZpV2
Ndv7ho0wHAkpKLZY960rXmpNfq6EN1BLJiN2M4usBdccSyiBdykUgM/KzHOlcdJOV9VUcxyV1c8j
STRg0UNNMhal/RXWqLeGHC7Cwok8AlPrEUmCoxq3nrD66lzixDWPcRtZDnnzkV+YdQNhYIIdLySU
Vln3kgxNDyf02LvUK2iqBi1oDooUloypNWsAYTVxGOp48N0u0zNMhUlxJuhgEIF+Bthqe6lYmdMK
rtB50JbjmycM09+01cu+ZKokcZeGAr7IUQVxzBA1ZxSUiP4SQkHhhYYNgIgocAs/+e656eMzWYC7
qsAhFI4JGfghjhz0SQE62hM7IN8Kg+qK0L3ccdI/LTRxwh/XNVZS3Xb1cGotYLwbjPPcIX86v4jr
p39c8LLItVvML7zi8mxF10C41ntXEupFTZRb562aThdRKRz57QHiJ1PeMSiPZnexpCVu8JeU1DpA
QKFt1Wzk9et8u+q3Nr5lPO597W5jp5tlE6U5kZl4uZZNTP3FCabSPkiEDTerxYVeCJRLLTOjNfbx
rQr36IaMFxIQrqHK4rUVzE0Vp2943FyVmYwKKb0yHaM3HIPYx5VSGZe0TbqhhVmWkmoAphu7Kx+N
ZNxFBXzYAxj/4oetc7FN/E47WT4paqgznL+weJMEPnOQgxkoYoLjwlkgLVRuD7VCWnTr2gElahLC
yJJpgRE+36Jrg9LzW9aikn6pQ43zXTErwRAfwQAMLUE5cvzsEfl4fzwPyasTpdT+rFygLn6mu9sQ
m3sDaBPGaqwGOuszdSFWGZFcAd0kH8N9lGW6rk65ekFRjUEuYU4u9rUB8LRuyUxxqOyNah73tkxJ
Vd0AE25PtuJHJbSDFBEmthMCzDT0D8T53Bor/j+p975RYaMx/DbLGUIRc+wlzubrgzaSm5BwL4kP
7WCGylQcTlRWm73ddm1fprXPbVp6t17zIpYrqgPwbHUSknFgCJSPoJXJWTjzb+Z1icIT2fRMKVXc
29RIYKYhZYOzUkNxf3Ek73UUdgnY//yuaEfSk3WCEOTPBUV7YN+bNEoTsd/zGSJOo3F05w71kU1T
H1qYIYGEPrPGa5LTi0Kq7s8UVqztdEOIc1Nd4oxiAmN9ccIe4i//YxyITRHmb/3jXH+dbs528rSa
8jqYOQ/Z27c9/2x1+A2PCp/Pe9wTvYxKuKCF1Wt5avyYs1Ve/DjFNzpB60N9R8EuvOE7VL4SfLE7
qATiOqquppleCELtc36utr7uSrVssJqQfzXv3nStnrCUfck7sSaOi0GVCGeUUZWdFcifqjoMao+C
AMHzyd6Sr0H9tleNY1L/Wmmk29/nJPkxbue6GmOAbUONZJr6mFWH6XOFHviioPUJ+mZLCusaID9l
7fH2aAvjBJZLhLdC7R6q2PqVJEikZIbUUjhv5GwEx4NItZDwNHiMohCyxtfalBwv+vmMtYaQPBJe
3vCLQ3FHeT8Io2HRXugaNzYcrzwC3de1sBpkKc0Xzvjj0lpKVVMnUE4bY8IAkZJpGQpzQCvfcdkf
5o+TCBtzaY5SYAJxZITgCduhBdxoYe1igLmJp1GVjuypRKw+LLokPCYFOUA6uuTSFm3A1bxO9nPp
OXXPPGPVq1HXkq5LXsyaZrDKyBI5RzvQPCRhsdV9VhvAtw35DoZ1SiUPms/zMhh6McnJLHadoGkJ
QSNlCQhPt5EiwFFfWvnLvzbDJAANjrjJh6dkbDkxT2tClwTkorH8H7D5+mPoaZppyav2zAE6y0l/
AMoSOYC0WPw6yG4WXLxbEHnOsKulf2xqES9mkcNtzwo8biv+SaLoYP14kFbqi6SLzT9JpfdlCtUR
RMkBfQBG/qW+FrzvOrtkFXLhKgfFWndxQuzroVFO2IdN33MonHQShOU5WJmQK0Vc3LvyFuwS1y0V
LVggz4X7c5IZY0aGTl6w0ptaeyNL+56ksHo3qXh3xG5Kw1gyZB5eGn+k3PYtTLsJJMMrpvLpzJYG
HkXRyxrtbhdLTzx+B6ihMZNJvl5q27Xh9Q5A503VjC8PhH/3tT4+v3CRu7QanOKzngpv9suXX8T4
tgMLKHADGllvFGMlQld8cI98UQNnEdCtHlhXyzAZEChh5ZJIi/aKJYlBy+dli0BFFi2GEc71P5M2
tzVmUfpiYfIpKS+adyit6IO5uYhhdgWKLFIm0AKvMj6veCVr/1HLghXOFcCe33SB0pZ9653aQAKi
NM6FWW0JrP/HJfmDJZ8LijmX/MUg2+meDNBdrKuKi027Wn3YhLmec/8ghgtUODFsbOtNS0JMITbM
wNcDEJRIaD1oTwV6SK8cB0p8+s43aPJ7gZdELZvRNrMkzPcdndxIwl8ZR8zktyfVm+FkIVYqsTtQ
+SomI2Ro2tKl8w0XUf6eM9v/6xhcyqkQCPfYxAXZgp7AcRR4YjJ6D536Q3GHNbuJ6rd0nAK/laSc
qNRuI/zdHJxvnqgbhF3UyOKtKJBZQlzw+kvezysgitN2Nt03X9M7YLIWS+HI+Py8V1wpZdRZRHyJ
2/MUG2I1g5U2PfShg/0=
`pragma protect end_protected
