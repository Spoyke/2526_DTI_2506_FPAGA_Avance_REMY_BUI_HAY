// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kru50cBE8uSSnAxky2K2G/ZJJAueDUycAlSmqBuXiaGS1qmV0+OT5UsM/Vl4BMEFyl5fOiav7YRT
+3CaQky+/reti42J6IGCDZ+cPhF9zt8Rr7w5v/WfxYiZ4FhMjDBidkDKaVdijtlYfO2t5j7NkdN/
N6eXLxiob+nPFDTApFHAuefoqv4QdSu7P/i+z4czcSPoXnkC5pQ95IU+LB3G5AW3gY4HeZv0coDG
vuUI9Op6dTN7W82TmpHym3EJnlM1QR2hSpFEQsoxTKpZ2qi69bmqQoKvQMshuFdSQUZmBm3MNyIc
2BVoOUvXOFJzNO4NWV01Nu7mVHi3om+4rkSUag==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 53728)
+zQmRCWFgrIEgJbuQaDUr9UKd0MQAO+ke0t4/dEp3cAOPPT7FLYdB+XGZ4iVSvvIbxhhzgsQdxIJ
yLr0sPCfgYUSUVm7oypQajM5tENG1cda4pid2+yF/h5KxI5/kHkdiCtt+J7Wwt29pVzKxdINcj3Z
KEHzRIWz5rTn2pBOpegCwK1ont2dQ7cvZ2UM1gxN9Okao0eGbqaY5ApwQ9+gibVZKSG78aqyiOfs
5HIpAKsbv0ULucbA7imUgnveLKJx3cxFdSTSBqhiqKJM8andLEW2dwt9iwSmIsRzfS88aIb8rbTW
OormyyVb2zJwsuEJWr6hjLDI5teJUzflsQJQyNDXjhcj2Gls0QCnyvDA1e1OT23Cd7HxMqMJK0Cf
1pKmHetNoHQ/ywaLc8n2f6OLZtVff+c4FDFlg8i7AkhLGqscoeP/LuvY3RN1yKeOtKeYoL3qG1eb
mSMX4lvlVDgw4owsn4rKlSqCZS6mQq/P3Dwx8k8rVlxVJJ1HNgppHQcDS7TFTPsYjFT2uqG2gnBL
ml2fUhLAISO8zC7CxrqKD1ymHAY/+llP6/ugOrJVTkwk/iSvAJrPsDFUADnwkk1LyelpFLb9gEUH
O5PW93r+IsO+xFOsHgG7MFTifr/uDgPaU5R5j6YUwtNflMxrqEUc8LZ8kgFUn5fY8M//2QUGr7MY
hCkSBL0SVf7xdTvfpIMZ3Np9eLrkbZKWgUap3Rpl9krOETQA66HMs033a+49qp3xZ7qnKXAkmYHF
9Zp+9MpfIO5K/m7Yu3yy+eAYnVOxRaxT9N3jcHvlVIQ5pOuVSQ4cvL43Q2qTcz6zE2WIhnOvfBdt
nOc/q44d8GyYiBMCf0Yl8nBOFeJUc2F4ZDimZ1Gs+8K/8brZS+YkksN/ZPjSHsuovYtI10Deznc9
K52bQTlozRdv6/im1WP65rJXplFYnW6DWfS9SGA+kvwhRDW4BE3l+baLJC1tEwQlUZUdn0fKdGzj
XET1jUQRU6C9FNBdaOTTtujQ7UU0gGdf01tJGqD8uK0wAEGciauodmwz6SMFxtokb+jGS6nAO0tN
YP26+Pp8shkC6Mh8x5ONDDe5iCKemE9US7ws8Ch9CwUmDI/eOy8dnk0kRPh5rJPaSgvFgzRDYPxi
s/sSkLNKXhgyAkDbiqHPakymS1TpxMRBOwiE1AqR8IHa/1/4a4YkADjCy4krrro7/XYnVUAwwwMV
+vG+IjTylqQu1TbpPMoi8imBOmVW+r4+e03S2gKaGMaCdEvW1nyWCQTAeSRHVAecaAc4dyC0HwYm
5NdjDFoThcOQ/sTAH3o4EoEYNVyIVfVS0X8Ui0YT7N0gBBd4LEAhVN/dyY3MijXzXnfzOFgLF9kA
Xn50SbUXN/IJRfj1WL5od6YiJJl3s/Smbsic6JSMR51ocG89yO062mKb7KVbiuAo4b8C9YDvOxxC
qouIuIO9XTSPXYMDn3yidIKkr0YgYfZbPevPnDWnnC65+buEgo7yXtPLecNlD2SVDvSIEzN4M5cm
c6sLUgtKRi2rPWENgBcT+Z7GMiCsEk2nPFMufH92HSpAGixNnAHel0PEhm3i5fuJGHvEwgbSho6G
myPRdhFwuksQJd1aGeA80STXbxW3bHcYc4CkFiKX3i5M706HXxy3/Kb49DTwgAqpNgxOu7rlU7tf
LRdEn6zCjFt/ivSX8aHNcOGYU6//syEQvQJ+VoKUkjtazaTTMT68dIVw7VhzTocJXotnUR3bmqau
4f53I7GqRsTTSM1/cst0m7lLydPrMdF3zkm0OY9tX06rxd0cBPcIfI5ZMtuQI6tj60r+NYmIXVsx
PrEjEE81X5nB9V/ysxBYblWuhnRvMHIWYNm9wbXyC+0MJGWI6zMueu7YKFNGJB70rNHul3yUgXM6
yQvL9lbw594Qtn3LCYIEUmH2TO3Q33uIrI9qqf0jQgcQ26bCWtcy4FEQ54vXuGTqi4zGGPJsvYDK
JHe/a1lq6BpIw+zot672dUf14yZRdfa3EWjQp+0+SCD/wJWPWLV0zkiUa0i4T5yfhFml5mMTVssQ
mvQ66xhzfQ8H3ybeEGbJlVr7Xvdt8Wgcr7o7Wb2jjnqAEce3thASgkno0eSp6/ON9O0aOmDmvyfQ
lAPZtkxaqUCb/lDUG0qwgMC8CSrtuyNA6gcSCqpHNsw6gOL+MsdEIpoQNvsZDS5b/dhrmaXzukEi
KEu6FLtZHHw+1KFyj0ydcC64qwoUMKTZE1cLTmCUnCBuKogGXZQjh0iR8HAJ4g6/I2BRdo4of6TZ
Z+DBc7Dy1GajlxTaV+s9hxF8zlAiXVkCu3ifaakpfjEgMJMUmwrmcdK0uqNYXZHj/fbOamGVtwbq
0sDM3GOumb0SbHnbul4O2igp4ChQwU16V9Agc8q/EGMxFMWcIf0zkdhApWHAIRNGo0wCP/JcyeJb
vQ+TDdatwuPyZDOxsKQ508JGi84NlaReBmBaZJVBv9u1OHjfDnf36ZHZsnezhlHUSZ8RKxkS/uRZ
MNoTqDgsyb1+6OxTCiv3k5VTh4+O2bo5fGRkCuyE+0VMK8nvpX4H/3kR+tA73o6BxPHa1ARvEtYp
L22S80QsCSt5I+O6yCxw4NEH+IED6zQ/ucHJiL9WBZX5yH9iAkC+2y9ZAGl67esI4tho/2F4MHH4
AXPuhj2bT7nRhAmHjLyEG6pZbMzkPdX1BnAkr7iRp+lTgn5cpkDPNK4GO3SjIxu+MdRcvi5pHqpw
HOG9dPeGsTTQHbYCgxVE7GaorxshFpA+41RVbGc9X8QIVMeE1cJBZCtXPtHDIR8dBvp6i3+gOj/K
WtxkkF6JDnw+MI+mZwLbWdHChoyk3f0oVKt5FI0pTQ2MbZ/JeWFH8k9Fm3mfFJhLDB2EsM5RDP8g
NmmNmPBzys/LGePEEU+UF4WErdBvaGIcAikVQwRESQZD5Ylp4//yjsE2Uux0EYwhJ1jy/pbXK/Eh
ClQfMxkAuEYELAvlD6tPIbTOzVvnwBxRUy8PFD2QHCtzgMWWctbDiiuHXiHUAlaIYaX+jjkm0pz8
w9m99eMt2JbYAQllHScJeAosVgjmZNyyviThtFYcXNJjFLI/Dg6DjZ7Wk2qb68hcaA19WFfuayZM
JyP8L6GeaGjft3k1KuTyTCpHWdX9aoPECGVlSr8QXahRmCCtxF++29CLtIelUueeMYJjuMJm0Syv
86DN3v6r3fYhQ+hIeHuI4yHxwXUUzasBhb8Lzqmbk2NzYPqV9nPyaj4rh5EFXZv5emDVUufpOdtq
MPL29EXJxTSUQ1G6M2PPc0Fjy7jzzl9bwH2GIc3DC7rbqoiZKqEPAjo2GE2wmzY/7i1xOBHWQwrv
baeoWMYhAG33XISPM/ycy0UIB2LnXzZ1TCj7ebfUVOk7xg4nnzZh2WXXJ5p2ZOKdsRSFw2GBvfva
FD+bZtou6kyMt46dHUvHTewdw9fuVdEDFDLUDjWS9FGsHaggr8InzYZBE5d5y+uS+QykRLQylPex
fHo68BBdNjTS5VXb8RNxNbOS6IGJ6ST1q4/lCP9ZfJhUNy+94Hx8A09aASi3aRm2VgVK52eCoipC
sSQcAM6jZ11dJUfpP/Pax6o1V8YXeLdz6ky9JrgGhwDuZTSXpj5u25faN7LuAJHsMTV1R6Wy6qyN
5tcopw40WWBz+MChElleAnA2K+74skGBrwGoVMumf1aOsC0Os194+6jtN6acD8477CU7VEPqa09H
wCrLae+lM5qeTZZdSa5QisDJnYKJpQbxjDN4ev9rWfH9ElsVOkvA91KbhFE3nxV5mgHjcHuZ0rKK
d1eJXWq7NZvo8Fa9sdLYnH9pqcFuSuPrgZDqMZ3eI1E/a7CsGB/MCHxK8WdR4kZYkrLpVF10yB0k
1zbLJ7wps0j9p+Wgr/YVe4ysdpYvpoE6W90OcS8SaLpK1SIQnRYcIlWN4N1Zm0hU7cS5NgLj/WA0
yVjbyUQU91gGMGGD6b2HU8H2Qv+9peJlU40eZp36nkde6X+hdxTX1V8RXFnKUBWqaR6BfrJC77Xz
x/WBaRMhLP2+fnMn2rOyzBcD9nLWGIR0FbPPYtYSnKHEMHJsAzU9j7KVwjQ3nCVTdBj9g0+nUBFR
837CdN+V3+5fSQLTfy935lrYTwBKfYBHhS0Ok24rneAjIu5/zy93gVd+8WOCUJXrZ+72i2ecGOgw
8eVOwUfaoWJPAmeN5PcoXuA6UrZySdSJg5yfplZ+61wGxlU++o2T+Pk97JJiq5Ezdg8mremCpRbP
Mtm9D5tKMMrAbHZjJb0GxpvZy26OCG6z9tqOsnIjiK2k1f576LHMCIeskuyNo91goTywHQLWcNBz
9VF+CAK3IWYvYqdHIT8mhaqX93JejlFZUsKrPjo/Thup7zLoTmjR3VBo6FXL7YP9kNU/ZecZTzej
xnvXaWCIfCe8Rfeo60gOv5HsmAJdBr8geZ20JV9OpvRjcC+0dHu1h3jg30EyB6YAx3hNpuYLnuT7
xLNM3CHO0gA5SMtfiX3JIpqzh1YPCbzDHjZuCF3sC28x34mK3bUT/TCZtzVAQBGx1tPG11V0xc5V
DTTZc7zLyKtUTRm4+nqLOkYuwYrWo7TLLrNZuccwRfDauQbRZCBJsUU/A76w6e2EVK720xpoabaH
Dpiz7gbk0dRqX1aek5w8xUvbcX9mYxTggC3WYHIgEU4bsWzB1ArBGm48KhJcKbfikaB2RUw27q0G
tAXlGT0Sgjxns9tuaNwQxDhG1hfy8sXnm69jejCEprYSMS29pZperjp9gGKcasz0r8LELNI8Oz6D
i3E5i9wBpvlP+CY0LAZvMz3PSmmRFFyusFET3egEKCZjcnHpQglvlz573eGZuugrJjITK3unSvOh
JNgPdejhX/okjxIySkrA6wRrd3vkDz4viBCi3Ak7YHiM0UUo0rgpionEZDyPLTc+Fo4CsFDXUiQH
GH+uOEyfPIKWFg3j086Zu0yZWDptL6VgONYsh62t6944RBrVRWLunK8qrqgvv8Mh1lXZVAY6F4id
gc9D1f67sNyEeWzWRH1g6xxYhFeMF4wKHJ/syVaF81Re8JOf1grnQvZQ0ukghkhRrD3GrKt570qN
AYErxyR4jqM5I1y5Shi8CtvsRljOqIbgrJhMqMEzrBxSoiU16m0vlHWJd3RpjwqMTrzAKxOOVoNW
ZpE3qH6lZanuHqgJvVxRo0gQME3FqFLhAv8v+BZWUeYmcZgRed5aKuaZ/GtixpTgto5hf8vjM3J+
jnC8ftk084DaepYggF3THYVOzv0VvKZKkI/49R6FjUQ+Rq5C/OEOIteXEP0xGhmvEFcQiYUFjjVt
bkIVczMdDeJ9labAWyN1Wwhj7ruJyZEZ71gj4G1DZOs1Y1Qdk2tpZ04P9k4L0fG4236xhoIdnsJ3
7IGCGGVxWLRMvpsLk0GYl9gso5yttWGDvnj4q5XbvwW4J9h1NXBNaKY4pjIbmmP3KJfGugX1pQDV
90MeziLRuDxr9hQVcWNmgWmrhTnG3XhsvfvOrF2ZqFoMDhA0liuhOaH65gYxewOXIQ5ziv5sw87I
+i2B9DIusRiwIZhIGXN//8Ih5IwJJ+eGLLazjmOjvy+Bacq7ghPxLxm6nACf9ITALDMqSoZstP8X
igEHna6pamBdsNlvIDptSbK5l+QfbB5cglfinAmBv89RXpXu3Ugl7QAUXSZdufpqSc57mBHSvlr4
/9K9K5GBhuVTNbr/Cb+3wk4x3FCFXlUZwJyuRPPCTIG+yCKO9/U3MW6vC8/IWdORANpL4tm4gR1p
THSqthPrLP2pE87ZadZEJoccJjujQbDEaJXfV6huHzZ3BuvE3TJp4Kc58gPmphetgO4TJb5/aI8c
uxX6Y7/eyIGG8tman1OWr8Kd37hvVlMQm/QGtl7BzPBsrQUKwpLK7lFhMzEX+GEmOlbmoE413q+N
kI8v5z6q9MhCBQfQ30p711yq6JxfywvjkAETMnEb50+MjEKgoIx/hS+z9I352cZp5u8AubkeQmC8
DEe61CGljpe3GnWE6VyCvT/uWwjrGSXE0jjstvCFhgShYDPb55TZsBsOmwkym854NaZcKFODNQCh
xU0qJxKEr1L7P/+P0iPbqQ520Drx2SxoKqJObvYoSRCbLLU8GXGDtkl1e50AHenWdI4KVsJOTE0J
RdNIOOGZ8OxLVbQMTgQAEpzhkoI/fG2e9YUGr2ugaUrqK3Ia5b3vQLhGBJ3rttGyHPxRvt7RtxYN
4g25hc9CuZDlt4rzo8WQFqmEEk0zVGw0xgioVZ88xfqdq63Nuf/ym9aMXuq+dUbJikn+zj7LU5HM
dDpl10oIxUGmaFmzdUGiQDPWkuVxnlwkdgCn0ISvZg0M/5n1txDxtXcIxXOX00QphjiRJoffbDg5
CGiXAbKEx0AsMpHC9mAorXPmjA+GseGequLW2r+zchqbdntjFXNusbfvRacZEC114ZupMwZ9vs8g
RTxboKnSy4DiIIYjaxrzPp7+G57NSSci6iPoW0kJsOTnVEpvfut6HnI3u37S1vFq0RX75xgjaiQU
AFaJXLKPUmklFg7aTIkql6MUG0OMwBUR3lt0kEiGPETTuC/fe6tiUHwMTc/dX4oGOQuRlWWgObwx
p6Ouh6gwhKciTg26IdGETFVIyWO2v9dt4JDCde0wtJvCH8eg99z6tluwFDxKlfgng2Es05deNABJ
JOaLIFyHeL6GgACjyBP2FROZSgKBVpBv22Tp19TiLtQOtkF09aUYp0EUUKgk0brlWGwULWYMQYfw
2ZoIUK0h2bJir5ibQgzgDmmC7+NkMCx8N6srcw8/axQSSYDx5sr8OwLgFBoTF8YWHnw5S5J13pu3
jzka+vaKZV51ACkD+VAEjHFIVF6ivIJlAuLBOG+vbJshYYH4QYAWn39x74+aFCzfPY3LZ1YDw7fQ
+7wssiCmnU19m2exy/h0DZIOEtSZVaBPtcCKGOb0Y7mICFUJJWFqxkuWvew3Go1MEqAIoxohuxej
mg/Yd3MRg2qdmgrbYbJsZbpgDhuYLOy6TqTEU/Tl6HiBo3tUMjoqA0qORRJ0eJZ4MsaGeh79LZhb
fxFn/BM9SWOVUfKWIjlrvgke1qlw6zdwzqTXWuEcXzM/TAZmGuet55k08r/rLsWIckNEqJss3zRU
cBN83ZS5yoy230lMpehoILXEbY3kK0QnhoIhwA1X7/RSHdHH0Y7Niyo0atXssqgJOaR40kUgcFCf
XDraOeqYlxkIZmqEEc10PTiTIUjSiQD3aJt79BnsoGf3SUiAFWQcMFvhPxd0i0lh72M8WtC4MB6U
JL0O8z+kanYBhP/3YIx1XiBoXEOFQUCh+7pJXcfs2XAkJUsPgccI0nFptwVT0sfal8nnJI10FyC/
hDLXxgLEFkPBxSbjagH2Jc3VCB+Or8UKf/U797O1rk3CM3OnPkcY4qaB4j+cGgmUNqK36MShYSSt
nCa4Z+8VRgwGWSsYdgaSIaEKts3R6qd267OGfMyYla+1Tw/50OddF0nutBqsdNx1uCqyI6W60jdJ
EGAwFjz7Bn56X88uIrD24zdqkwcX7HUAegcUTiJC/8PxJx7WeA0CE1g0EU+OzcfScuM96+5NCFLT
Xq1TDr56W8qLK5m4Jho0EBEsniBSn4gDpA93wIL1dLLl5VD7eRi+6CT2oBMN/F5vFP6fa4jyLM+S
4W2idGelHOmZxrxcGijm1+igzEconJocHLDn6VQMPc6cJISVDt7Fw80t+vimqxncwjB5qDO1UZxN
8hrBZNEq1Pw5FAWZtjoC5JI+Wy52kMbFYbAsExrtSuE1cFXNhYpdUqqQvtgE0d5aLMt0P9CuleCK
TFmpSHMp8HR0AIn3rYGkkZ2PJdLicT6oD5Un18ODTscqfKuKHkkQ0PSVhMIY8bpt5srpZE8i55/C
g8QD1idG4sEfiUkwxEdpraO69mLDkzl80RmuGWg/8dKGCS9qowc19jFxKBXcD1hTgL6T841WrN3A
8v5K/YhlqzD2pp/vctjhvpsfY8LltAAFPFxJ0WUF19FuQlaYPSzJ+yvQpXXtwtKXkSujzp+dug7p
oq4vQvmfAnp4FaM2LqmURJiFE+aZia5V7PEkqRzrlSmiEh+0V8sELBqb2W77Py0Fu/dOptqPXJaf
GKzRUSd7t450uvGeRE2cQZHQNeVPEBZL/4URMTETPE4uYDIh/egGGgrStShzr5O8m86EpQU7dPGj
VPgEizouBHi4pbdZXMCeD3J0T4IIa3bgjj606rZbjL1TVyOX32sOdvI5YVtBLZjJRcD9yTt+nBJZ
DPyRwDFvGaUkGFxxVI0hjkWzSWCd6JomAUN1M3ilcnWJJJtBrfP4D6+6UdhaOePQlvXtBg4L5hzJ
1Bq+/wItwl45Ts8OlqoaAjBH/bUKjcrk0uhUonGVOXXr+xdTDQCb1USTpgGmxu24Oto+RwIV81+t
QHb4FYAmaqy6PP+R4HSH/JMthd911qX3EV6hphVNxPh1ntBfVdjIVSCGnPVwdBOsKjzJRzMQzzmR
tA3vpEvttoXtjZLQZrXceH3njCkJbOhnKKDHh81WwTrkXFrwXuKCdY7XxAhaOnCdEJXWp2CjQ04A
WLnOqDp0RRy+d0f5R0xazfc8Q0VFUSzhhRgkI9cyrueOCsjMBC6pgQZtlObY09UvWJCeK54yOXPR
P3BDvYxTJLJ27jVVXQGBnRL4414Z/eIXTDF3SxSaXD00Wmbr0vbX8epapUWj7jzfRwvAhWfHfBxG
iyT8KnY62ZRRHkghZSqzMwKV7jXI8C/VIe8k64rx+Zo/b2ruTbTSW6mM95gsYPQFxbXBJUboSTTZ
8HKYkfi/IME6Rt8mvTP/eWMDTa9JO6D4H7u1keXT+tTnQeabcH0avwdKjpkRw5Qlt1wvPPblpjJA
Vn6AzN8ueEMbRLyiGSiOyzpufILCT3NpBuKx3N/4EjB3zrp2dUsZYTQIjSkwkv0E3MCH72tdwbTS
WnDIYqsBFt5O3u1AudZJMwzEE9FW/sAFsNYzyHyAGXuKAXXr6DBAHphJVUFHfAM0FPputV+5FvYV
ymRazSpolvo3va4FaX5yKfVRPy74RbVEoyqVDCjLQNlkzsbTk2NKegxUJyhSURvSOaUiF+WjKqok
zrGLE32X/teAt0QlqniK9oHUPi1tKXK83esKZI0WPdZlvM43k/sB43sSqDjBp8y6yKexBjpItQqy
HFhygch7ffqjXZyAE2qpKAcD4YP4D39ozybmhHJsist2TFhPHoyN98B1jQpUmrGkCeESab9MWL8I
rHQYb5VlGWx8e6HV4J+NshzfC/P0Zyb9bkAegoCUAgcs6EfI3yr1ENLSTTaVuACdOEBSMuwiUzjL
oYDTWRmvoAHTJvVOltwDztrwx9RA/O7kT9iBwgrqsOAdaRCUMnhRX+boJONYEoopUwB8G57WmVea
xOkchehqSbTQum6wWau9moVtzjTEsABAQgeAR5RsIQVWNrrcjTMzGh9IV1V8Ee5b1tR7Y6aU65PD
q8Zec2udM8sbXGI38x7BM7LooHq/fpMW1vCtfTLik8Rvu1fLSKld01eDtHzzHKLqdzlk60OGZ4hs
bAKU1vru/LjvFzSgVmrCDLMSKRDuUWDjnUlnfoCPQzhjcVLt61poYq/8CeZIpZSbi4CvRUVXZl1z
/iZJpxohLVqceEAo6B6J2gqRo3QQV9035mYIw4+dfeYew94ajBCiL3L+JpDUqjox/OcWBPQCkRqD
qJQgO4Goj0SEszlgXJmIaoH0ZrNFNEDpafrs2AQnfTU/dBBndG85sfLLLltqxXZ+CZFkYW4FbOI+
BOAMCWP7HgJosD0W1MFCpiyfZYkR/2bbN76UHSZHIW+R7sVfF1TS0Q8/30ly5IVcF45f5TO2/xhy
Xj218mSM39HpGo+V0KKJrkXYMqHM1f5Rb+idEZ8zQR8ThT75PK6LVaeTgCuTYVQQVBpbg4m1riJf
k5DtlQmqbhiJZxvUCeIUOw4tiwil2/bc8M79NaGvIffFVZ0FA01bjut5puNzvcINGBr7CGYcxg7F
uyHO3n5dU3zBF9uBf7Qwztd0VxrhoR0swsWgqNDLrrapwrxxpdyQIxEL3j0AV0jw1MrzU9ueOsgH
sPg9ZbYFLGreiakGWIJ4rEGgXL5oJqlARhaLWc+B0rRoN3FU+AWggX7wNOkMtLkqA6sWv3pqRMjT
NbZ9JN0cZXjk1lNMwia1RjJDCgwLM4J8pQVPUfATiOT4pO6slCO4yW27c7c01Va3IHO7H9VnjWNJ
vhgUyT132ecZPg6qm6iXQ5sKpK6iwP8aufMrJD4SX7IGlkFlZcNY0ELOPtpRZUxqZ9PyK010u8IL
v4qoSSOrHhvCYtbOVf570fA8i19tetggsrp0E+H0HIcimyzy4TzmJc6rPc/bsvVchIxrg529f5Ih
H/GsPMEDTAPUj9QaATPgBHKirbLsHNDCALRCKySZH6A8qijq39N0DCeQ29NRJaj4/P7SC9LricEY
J/X9PyFw2Ae9/ueZnKDPqQLXFkkEhUnkKdxNObPQy3nXLslV7sy9GZpMwxLhQgqbFplwJbgnoeZI
l3mGUgdz7hGOfrkGr13lAx6Qlch6wZ05CnlfqknPKo9qDmdT/tGcL8ZnGKOIc00mE7J57oqtHjus
3oG5XIh4GVBodq/U9E4385kkcTopyjdTF4w6t9ZQsUry4a2zmBnhYgRez+WNLPzfI+6zqF0jz2us
q/4WWMrNw1KzljzasZg5lQYZzLFEb2l71diCBX/UdMFjEYWTfts6Y400A9y24r9S+Y2yaCKxJRYF
M9qqzoW20CIvjZN13L+6KEBidqs+i3mkVdQRupxUWLMe3CENjRBULJj+ujFQiCQ7VG3T/g6Qv7Si
EecPDzvgfXgenHcP8LLvQUSTk8YgbcISmaQKdU2D+096Qefsf2dLMhlCGmGIdPUxFPdPrMa8WlxC
TJ9Tl9x5dbpN/OF8L1xnRaGSUKCWdl8TQiKIp0mi96qhUm08KJQ+hdVOa4iiwn56hLODN/pL0Te3
MaY5ygiU7VHUnYYTw7W4B1OY0GBx26r8Zgvl9h+xuUh3VqAmmiA/vPgJ3itMCQ0+/SrXlqZi+o9x
TAORycyCAU/on4LU4WgvDAUyCbH9yNXj+dvKfoO2MNleQta3D642oX/yvc8X+7/1WkbBdQjoap5X
imwmqPhT6pxoTTl64yrDidgikHUD42Ocgy0ctAHjVPR0U4bGbNDXOveVpfvphjK4SRT009w5fV09
KgT70u3ujWsbSDBlxiDZfwSaVpPfc4d/xEXhnkYUO5uhBvqv0qwo2q6r/P08y3nFtxK7NDox1joQ
ajxXalNMz7A4/oyoDNrzSE1HwBopuxKGKcEmW87vwugFG9vaGCbqlvgzY1QXlVjUFjB18P2Z4sED
/H9nTQOuqvGkhaZIsGYbRmvCFfNf+VrkXzKbtAFn5rkSeyfPhDXGZzGrelXAGjabck3PkpvC2i4L
CMgknPQzd75UQHISuLoVuu7ar1TDMCpGvgpnTmfK+kXHtSZctPZKm/wfQ+wEEPT995ddQtR25c+Q
bcvwS1+Y+XNpGvCl1Ru2NfWVYf6qoFb8E+JyDcNY8yE+ig518nbl3Wzhhjs3lL0BYFJh9H6rZxvY
0kgSM6lCRniPUKrL2+fTdkKfmwG6Ej3dACwYa2SFzNknaT7Bu+xynFUadqUKrw1uDsG4IlZse7Sq
+kFVft+B0SnoupS6uLsr4NceMDY3DHDHDlbCQFi47M4gyY34w8uT5uEEliSUk9WZ2PnYEmXjRLfc
N23ADKsEwNHGDPYPFWrv9un2MMLJ5P2xt9rRpMW4hoHTze+DgM88sx7tQ7zeDD5ljQwIxj0OKYK+
gEHCNYIvWOKX4S8nawax/PRP4t44wE9JteZhP3RRs3WfPhjVKQaAFPYPi9VoPgixCnObdruky5z6
770U2X96Q5gB1wcexQX02smgLnU/SO6NUZVT7DG2+8WdoiXLIQtgPZDyNLsMhnQ3K6IHbc9GTU3C
oLygZmZh9/Tt3iUk3jj82CteNw5vfGsvs1EPSutIIBexBQjWg14/buCSZmHyGwjm9w6T0oSrs6iz
KXM4VNDgJReLHWuelyQmBEvE4cE3eTaEr2UeeQ97iuxFG9QsnXu8pS+UPMbwu8jXBVaE+3D0wFME
o4NrQZblCzeAD0l6TIbo0Hu0pzB9LvW5IL4iIS28HSwlGdIryGTDuyIppe5aiFZ1vN6eGyK2lfvM
q0Uqsrg8w1+3OYPjkTfLGVR4JUFrNExE3+iwM8JLQhsonJzo60wSrdjzj7vbkt68Zabp+x2GNZwn
j+BlgbA4mz40Y6IoNCvfWnttl8mtRsXOo5Oni1yrrMRxfOQdmI0ugKJOB/XXBimxEqeWu2fK2dyr
mk2EzT42LD1p0Cg5CnAthSwkkYmNDVXEwlNxYT3y9R0UITnzG5co+eoB1uVXB6pzEcHAjRTOG5oG
NlR8VX/QJj4ockOpwcIanqN38kWVYG8NFGWdnMnKD78e5ZPVdsiEHms709Z7AA1XXfIvCbqxpz7x
8Ubl4DqowHOvyiEvYbxOz90mUn3iRBgH8BdSzgvtvKs88LVqdbaZqVpnSMAnNLVc/L6g51M2jZQ2
UNUpHEggET0geW985tZuyXC94w3ltwbyBuO7eqeFbHDJ2UtXznFkxudv7d9FCsOF+lyrdmfEivx5
rQu1DC1sgqmJ/qWqADXCJBprmasBDQUKCytkQJFvKqT8OpiBmfSSJpvczZh8VHqvwa0dCk9+MBVi
WK05UmAZm4Uq+k8O6LB++yLi8oByBtWWvep9LDcIFmSXFd7hyjR59L/INUT1HXiMwZD4eKAjBAp9
iF150TYOlLQ7Q/m/SOgCPFG4b7ZZO5HVjhWm5wVEqgQMSxXKFlIbvVdttlDRgz8JhYccG0IbQDWf
h9OdUewpjtmy/kHz6bTSOYF8PMFtlEFUvA6C2NyKzsd6x/PkxqprxD2IebzRoMF+pD76yJOMhfq/
zYnYfwOnY9TTyhaALhPedV7k0sRolwsYudqWSj0ML8alkHCmZyGRpbMQtOpBC3F13A3lGPa/qR2a
RX8vNw3SP6f+0BWsY3RnfTCWt2DAMg4NyNhxujLsI0PFteHNascF3jM8acdF5+ljwBfJ+zRJeld/
djXv142oM99i2oNFBd+JCGDv8ukdfcc854CWfqy3TLlxpC0yNQgPPU2JngfixsfBPHjAjSqwrwi3
3jY4D+zvDWNrJzI/FQqI6MR2kzJ3V5wgAqzYGgdfuPLFx+kJvf+QbLx2NQ4XkekYozr499S3IAqX
EU3UkARPFqKAX3ydw2fpodV8AWz06mXBpQly+5OOSGGbPxt925NrDj3JcAxz6+D+F5KKKvfPgIZa
7Vrrevze8DGKd+HWrvVV8GSVBFcXZZWmxchMbwTuYgsLPXDHd/TBUsVIXNIKf4/Zh2mNqStGwWsR
jieOS57l3q7ISnbprerdmWR1gWVdJ3Aogtx96Y3dhFTGNbPM4OA2K1gJP2Wb6p8JNIGYZIrB8fLw
K1zt/HIP/mTX1y2YRahmz5A95s+MRjwS0iHnLhnK4LY6LqV2Uqv2OZCDU7qVLgaayarSX/fMwKOt
IizFD7d52xQKCi0b6gz5YHd5YiLkbEwgF8E2eWO15+C9h+0qnVbvVXxfSovH2i3dfYJo6y5gV2gP
wbiHg5dAfmOpO7qj3KYOBddl7mxr0y3OaA7P/vsUPgWwLWKEqZMt0Yv1d3ctRxeGeNFfMWIis68G
vkgppexWku6mkthceJDcrpCHeQQu6a3ctCHVj6qm4hUSUjTfJKhBhsB9xfy3QvUqn692+EPdXuuQ
iQ8sdmhCGcLfJ7cVoCR2torVlFJueog7VwcdBgkHknK8dXe/hecoqNeCBcBasdtWQIpu1kEHjXJl
YPSw8pvz65w4T+aw5/ERzE/OMdS+DCebGW3LeCjL1NjHQVdw22QjbGYto3gOYDVNh8VbwNF5+0oI
fOsNChggPFrsv8repat8nRztIclJgb6qoNrg6rXr1feoiLghptHZZS89mktyj+RCbA0vMfPLW4Xh
k4gJ9BAb///kL5yZPKzU0wv6ojoNPqA9rYErpv2s6weXAbpnFc58Kl+E4FZPiGh35k32GOTBBNWa
TqhXpoMtLiga5MZcQB+6n5evkusJa1lO+M/pDXX9Hjg1akJlBiegJYboHGYazlztkArK7zmUPU0Y
yTMh2PdTi4qksLP81Su52Sotx5abYFGTrxucF5LehLruAuXACWHRiXv0baOFEE5sRBhAqsccNkUA
z/CdRABn/yfX836Zp1LQWFOsVZWNvxE9iWPaHN9B1m1tY2ax2iuVZFKQk941xyMwqGSQuHdHVPw1
1IkHYkQWVQZEdL+pGdjrhhQBADFO6ogKtspN+kuAWQOZbMrmRzCAgM3NSe+44USVxpB9CVGW9jg+
PLdOyA546s9h0YlLo3e4eNr+AtvLNcKu7MZzyofzkPyq1kZv5JTAR9CBkFNoj1LFyddnA22IkHQR
3zxScrPn5V+4XogFCwRIWxeUe930cIt+TaMOq6XS5nZotUUWUB2AluiJOStYkO8IhoBrt7leF9nW
GJw505+2J3lZq1aaoKexlSqg9b9lNgFSHFHbAU+KOgWzAtrGfNHUuklRvdZoIY7la2T0+tPkhW2Y
UDts2kBG/49S5DhQiTjiZbJpz9+S1WAlUas4U4zMGscTuZ7L1ZnUxEzSnwES5hOq8ddn2SW+awMm
Th+FUeSPVOH4eLNOx2k7aCFo6xVE485WR1/ifOod3NZHrmBcU7g2U21kIuVfb33WF3HrLkSlGKwM
VbC7MAeqHcKYqcidarpiqrndTxYKu6VGjNHJg0GNaOdnwpQAIaCULs4c54ZRpejCXWOqxgPis24p
3CBKpahhjWAQl0zmQBRqNpNSweLKYBFQCk5VyIoukb576IE3hjkfBYol+v78bRtN0DytbuXGfkAY
0utT3lyIM5TuvF1WN9XgB3lLylUCcZgJfRAp9kE9UFRG8E06bHEk6XXhaMg/LDuGY1/Yql4dTVZm
vQ8bpgjjgxVKMAlwfHrJUSca8sGqBEEeok0bHBpYvdBdeNqfNm1Q0XyZngUrx+MGGi7wVgehDdKC
UMUfMpripRBwtdHsMEEMxxg+D2vUVjSjfdoUf3xSgbCOGCR7IbpFoaOZg+bqGyQbLqBLfJeISw2i
fEw812S1gjs5t9jmWx/Xuur2Tl+ZScl5y2PGijUKA6ZsWln03KRDq7jpoBgtB8BUJWNxz8ohdqFo
jYw5bWtw3yBowFrqECyVUyVfk/5LTRfkuZVPqClA99sej0n+Qcr49/uxME/BU+gvgdM7r+4biTiM
qDMfVmIVPMjzezCCFoiz77B75earnZuqRjvTA0NlnrMDJpJMIUCe9rKaWuXIX5WLKfC6S7J60h2V
hgmZsdNAAmoZ3dbPn0mm5slIqMDEE7VDdcAg+4/iYrVcaL3dW4Kf9+Jqx1shrWGNj7Twhmd+bDBp
yRaPy6+zNp3j4UqO630HRvZ/dqU5Boyg0hE5eomW9GT7rGnQ9asEuwNhtNgs6nvLPc/VlAnm1Tah
pnOh8OIL752BL019lE/nperzxr3ImfxM+7JsIMEZwUMkzuFYKfxlLOKe6/vvv+0xiyOx18/kPOJ0
NZ2e7p3SNo8TcNijje1C50WPstjdocMRe9z5ZYEsyndwF6DR8IzCOGAuly4nFV+kxybTrjrKxJu9
WKBekSwzxd88xfwhgby65mq6JqMFRtah1RK7TF9dRhsyQ+/Zh4BScobXwLmQzxjIsJKwLTrmfWy2
DW6VI1EX1RwGB236B/U2vw3o5xAgF2D5ZUO0t54AKpNiifFCL+6OTZnuC8HxcmVyN/qt0tAATIsZ
cJ0mdu+/L92nnKGfd7hL0HH6ixBG3vS4Z8gLKY9OTKq3EQ1KWlCxrnhSZGq+Wn5ppJvS/I0x/uXF
8B/gsTbnpWjMNIgdSrc7EtVwd6GXERFDgykaWIMZU2vKNhmnHRlr93FOHb2MjfRrIiW/9AqbrXrJ
URMy6yNSGnIIgjLwKxelYCIvulawRXT1qy+79msG4N+uqXyVgp4ExfPy0IIwhOpwmhfH784p2mXP
RGiGZLRSyD+gpAngQq1ODMNzgb6jAJ+6wIA+hM85g/NMiNVmgqJ8SHeMRzGLFIrYfvBrL0q715cQ
s2CreG0KWSmag4uHR/R8eXg9gMERM6YgoQnBpa3wAaqwqpa551CdBqFAWvZvX2r4NnSozKJETzPL
PpfyJSYmYgfLvB72cYnLpFySLbfTW0gw8t8xtRS9ZHdmBQ+ifw2n5uw3yYBnmHiRRsDvUrnzx4Od
875RhX7tz/blH9HaJMo81ZVxhSxs2TLdCEA7iTGMSk1sDmOXXimet6AIWh36uDBPRY1mfJvzD+gM
JSxsBfcurN5y/HjRvn/s3Wh1cGJF+q/HD5cqk/Ui9qJgg7oo4IkvzV/DlNpKEhbpC6gZuhD3UlOk
tLmc+U0QFzak8hAQxhKMxzOFm0aMn5LJ/7yNF5SAJ/3hatxuOWgVPX8Zeo8GFsr9BCMAkb4ge5ks
jIdtwtYJXjkieais1gNDrm2g3lS5epAmrekO80c+blCGNI1ApoSB/GFqf93BTChLvfrDLSugM4N6
qvbI/NjKgWfWfdHN4u9flQSs/35O4ZTgxDi7HSD6UAIvsUL0Brnuhem4neYlWLoRLheM2l6xVmxk
7W7MZakGk4pvXU30Hr2TsbNJh6a4/3UjO9TXh1kcM58xwUeAqNrzVKq0yWzQF5u5J3IxxFqbymGi
zDTci04JsFTJ0llFO+VUiEUWwDNtV9cnFyMp00IBC2TEkjryTNWjXGe94CHX0xN11QYAe6ovTT6z
8ir9XW2Dm7VPGKFqpi2xWEt8ML3cogDhTOV1LKfYYonLIaYvLMUecQBENLE9+UCjXq7Wcy4ZrmWl
D+f2ZrfV83fo/Py3CzCbY5qYl89rj4JmZIskefvhCGN7QtFzI8po2b0tFtJ7jImPgFa/+TqpNMI2
cy1vrlClCOiQ+6hUKEsJ8K3++YtrcgiLa0rc2g2+EBmqmEV0SSZjjqfO2+GCo6yDumMWALBltvQ1
2Vz0fvMpMokP3ewPzSm4KPZNH1aovzQY7XqSWcQiUTCF42MqSwqG7KmVvLwaEIFEWDZXyc8PrrgJ
VONemYvo4eMoG69M0Jw9EwCO6nOgaGjiLSML6nSllFLQeGWFwYS9F0KMGr9M22JM5FpeXoQ+/DEe
6ApPaZnvG5oqkGwSL1XigR9sVafSpuJM+iKO3U7FjU+yspczN+/423BJHv5PWkqrv/8byvIGXYJS
kvIBCamlJfhbVKgttDGlTTHJG7IHde6O93wvvfrpXCIqtz7zIGoJvHlaP760Pxm4OlTYA2hb0tTn
FbNiJlUYdfJdrHt4QBPQm+RA/wviessRRAW7PW7fAektjgwvyZkvEWDRtBCR6xqh6arLcp7PBLY8
Lrn38yvu42AOma9dSN7Pwd8y+mtmVpSkUyyLrl3a28EHQ7s/8bSf+7hIlCc9tR0CAZYPrVoWEUv4
Gz9Dkdf3JqePhy9GWHhRPb8GeLiB3H3MxWfUK1iND+pLhCdxMg8GKwwxLAvRt+9fx2mXbZPyFe7b
PWKa/Q3uxBwCgGUBGG2xL+aK5cXqSH6Irg16hbg0XghcZRm3TflH2xy3S99TupZPp0j37Lfl7ter
hCqsS1if3oAAuMzHDhmgduhjIa5Cvu9pPRuWO6IDA/T1IAzqvD1toMgWlQQ+tw59n3y4r+oi+A4V
ISYT6V99Wjk75hPwchZvx9SURfhBqJ+C/3Ve6lfLDD/oO/o0BuKut3FJwNSoXKHArkCop04NNZlu
Z7OAbqso+ECzKZs6Ns2kmiFBNvCPWEGkNhSERTVF2l25jNeGe/uToLVwKsgE0Vm7KXft+9Hr3ZRF
QPpjlu1slaMrnXUy0kj4TJOWxHhpmUjiaHQ+02rnKaRSW3Tww+QXKW9GB7Tzea5dFaaT2e3xQMNT
lhbYfXMYd74d4vbI+XfRT9zjSBlin4nyrlldmHSC6OI0whZV+vubU48LV9XKx/mFzB3d2Wf7Y2Bf
tcC4LrIZuCV9f8MUi5FinUmvYoKSiEd6LAMLWfRZ0nYdVJjqd1lkH+e1TQVFLhq6TzR7+MIOpqdm
qskXwoXeMBYFCU9V3Q42egLNLf6p4JPIV2vD9XF/zd4JzoKssZeYiU/K6XGzGr9UHAemDCp9Hgmg
2uAjsYNfumBffO5JGWrxuOIrojCOv2v+Q9FYIQSOMzfUjdc+OUj3DdeLkG29jIO8nI2zJ5r372nB
vuB0xKu2JXQIsFDXWZw72fJq7o76Xx81tMLMwhmz1t4yg5O6G+IxedUsdD1ejaSHdxwbOxOKpN2E
N4qgjPHSy6n2Co94pRC58pcfC5p+GoOF696WpJGY5/d3RVA5Y3qDNPPN9cp06ROjvBgv65tbQjW0
dog2nwxGrKEl1v0ry5MlypeJ6fiJhWij6sFV+OOaEk5jvfEqfcGB72QPD0/eVhmkJkJm5xeTJB+n
usilY03I3CVM/2Jf8TVGBRDgfOigfjJ8NgPwD6/0lExmlLfkDfS5ldZlrq7J86DDltwZSzXn4LiD
GttHrLkHooJbCx9xF/VhpxqYi0JWlccufYr3Z1UfxAhvc3/XqR7/MGZvOQIcT9AnwFEAN2o+va06
mzVVEogl8LGsQMUj/uMfDWgiTJMCFZRepb3IYP9IFuJNv3vTmJ1OxmPqBT1cMyJBURKku/AZ+ryg
EnEsBg3fP571htvDoPgHwFmHK1XEKbbuXMk8r053unLerStH8+C1/8BAdXpMbZNDnLCTSKKF3DFi
EZJ9vUq67GcW/VTyxInG5gNVwjeaj8I1T7U/nOzQzOP6t/6rQlF2DlBtXd6Gh4hMfHk3uZwgTGzL
LWiTQuZL+fA84cq8U4f7Y9btDpc8x03HgZe+03N39BrMW3hP3dwTfTiFwMqNAo/+OQdA7Iob/bM5
UJNurqwVkrUyvLqdUT5/3SIaTWIApwc47XBCwsmzn5anmsF/D9D6q5hNw1azCim0whmiFfAYVqiB
FRzJGzBhk3CaA7UtO80qGn/6OUUZsNxF4ZYxscUaqC6rYw387zKo/uQHiZ46qsHuwmtnpDl/lA01
EkRPXoH7WWkWm7prRdwCLE0BBl7jYuRFaQl//DVasMWF6LWKW9ZStm/NyAawfHAUnCysfnD5/Ohv
Hy8buIhbUdWLzU02hrxmRW8Di9EFrzQjNy0yS5D02drCmBfrYO+zYc2fZQVoanTAZP9ATOwFO+Ih
ILb3s8963UvVX5cfuScxHl7x/5pOeC1HwFe+TlcP3bFy4ay4+8Zxeo/RUsm0ZM5LyfW4VluJPd9e
S9n36EKiLuGKWhHSG3dB5x4LRiJOrPxV7+OHNSuJiMWVKWI0rkC6AJwoR+Vi3t1j1jGjZvv//NcN
Q6qUDxdTYDdanmaXiPI2ttboeecfOUSV6C2H+RlppH6e9y9Xjx7+WKV7nUDflh6O0rKBdEQ5bLPl
nuYGeO6RDTJXKtxfrGm2DpiLVkYZk7g5itXJ0Ooi/yOHtMpazlEhvfa8zMJH+9vTE/4vyejcNurP
bic+aN+uIGgUuwTcxtdxYnM7ys8ehir2+gujpzlugv4cySyOR8kimkQXl0xJ30prdJeuNYyFOKma
tEjCzJ66HEidilh0GbzrxPUVhcjrEz9VAGS5Kr7nSRZ5UKTB0wQ8ypF1OyV3q6MGTfRJ+cQM+e7/
CFr9phdC+47F00Nsa8NVamwjxU42VhpDFTufAh+Mdze7FvNC8Wx3Lt7epTPXxpl5XsGSORek5tDV
UDV6GJeKnc2V5X2WFzq+kGIkY1HDHIANlB/BdB8noQr5wJRKdS1M9C1XHe2J5jwMbYVD0BywJExC
lt8eabrY+KJIHmuQX4fg5Vy+sed+Z9qSVBvU+/PlkrtIMUoALTndqZmBqwX5QLQ7n9/ngW6WUhzE
tu1PLoS03v6KkD4tacM2BBAaxIZtmXfVuYP4lJykIo0qR2ZSYjbLq5GjmvuZAv6+SKSOt3yVoYns
+X4f2i9jQJCHYI3KfxXwU96ED+eHHqdoZBTidnyDzcrAdBtVZ7OfVymDzJWGxyIGJMPjW68IfCnB
WBtA66Bx8gipDph36RmDC17EQU3+ie513qaz9D4pI3dUHfUB1vqjIBwgTG3zyPrzdZBYA+bqm15s
wy35rqtD+edvNKldQsrK2qC3crOnPri7Ch0koWfC/jUERmgWGM5jUNIa/mHn6iU/MULFpFkZb8gQ
C4VgdUcb/Cjpo5zALQ4UlSfYP1IMQyiGk5RlA7wR0hZoJMZazsNuECgAtYBuMe6+hn8t84o6z6TK
S5OVaMXBwjEFvYiIbG2/GYy65tcqCoT3LjGGp4PkMduHEGSXd6RcR2OHmDN37zmxRZUMFe0wrhYY
QWCmXoQNVaJ+S4ryrvomjNPKPwYMOysaSifrXV/6H8hcAX/njEdxHey+llPsQFmRDlq7bRrHe091
JA3XSKcrZbvnWPH5FW+rcfhLzX3gwIgSfpwsBVG7emhBTZ14c2xvsLLTleKtagwqiDJKxtR2KFuT
RvNEKOF2a882eedkHX5WqN6kXRrt+5c96zwmUQMc5fTeDOUMI2VqPT6GMfirNW8q8/6+5q+iIpz3
3tZFIs/v5J8Xnr9agN6QPqzWQZet2vZOCNwF8B3hOXMVzRreuisNxiZjmkQsNj52AVuqkwXJCFca
BHzHIlLFLhb8gOOvlHXdUTTVUZpCDreI2rCiXu9+EXwB58sL4Eu6qtqZ/TpKz0Me8T2pmF4w5u1q
HmB/kEkPAsTJdodi/q+WGc3xm+wuMNGM29ZS0z9F81uBkOfnNm0j9XJKeLjHyST4fRzaP/+5ifvt
5j0NUrb3T/MBuoB7bWZds4yG8LobObKc5sDQfuNwJ0sxT0BwP3PMFAWAR9BdrCOYJxNQYPgpsgFU
b1uTU6uHTaD3/jh7Mn1UpRvVheQvBf7xaLN7xyfxWcT9y74gCu97mJQy94eKV4PzY/XCRGMUkDnn
9zO7dEMe2Vy1/iqimm9RMCQuIe9db0q7L5b+q4eQpbl3qgd5g2577zxK0jQvVLma+woAtxuR0F7v
tXB25S05PrVqFIOSSqVd3oseUK99m7cSsdvG7sRc3Ij5UMjhb+6u0leHQaDU5waXED0GYFINRALg
LSNR/vbtQxxHIi/aTGdQYxMGb8BYqwFJvuHtzkAhZMvCLdvj1xSpdBVlfmFTkpCw2CFhxQKQb2L0
OusMKJC2Wvov6NawC3buLCJGkoKH0wNTNPDEMQNHQbVQGIDgyM8yJendHMvsRMRthuOVCUAzcBlP
5sK8f4PTXpWPKdQc/ioXO7o0/OfigEarp16XFZKkqoLeK7URO/3UEWalvEyBTSenAf2dpjOSt83A
5AsusWlltu+8JPXQlptZBNAeUpgvJJ9Zb+wWue3qOUUr4j/olpe8887hh2S/C9s55b8Sv0T2WPGn
WpAUeE0ObSCpVaj9VjIRfnLleUYNyJaClCJQgrQCN2VKyq3EWabVVsUUJvCqd3HTedt5Tb2GgOU1
UNrZNTpdmFy1z+lyNDeZmcSmuWNwMU1FSTZLuMZe5LhSe7kfz/+LspgL2xseKGy56RqHAX3RxNWd
yiF6SZFV6DA+bx2r/wW+uxabgdnhCtkkxSWvFeyZeEQ8Dd8RlVgB110HNBL3NCvX1yj1UaNfwxZw
zMahD6UCoEhg99lp++TRhyEWrWhzwPgqblm41BeI8eCk7e3z+7QXf8kAJFFLHQ7k/EAXmwfGIqrG
+zei5jHyiVTKLmSOCK1OlZzb4rnm5QRw2W5/NNiMj17c20YSXN6TUs9OvD6Od0CXy9S2D1bak4EC
+ppTbgnsl7JvNqt0OSrHdVpzgvuhi1HVpF4UhnL6f9vzcUwL1I0D+RfwG9/CyREMQTFZ5mSrawZp
ZXpHvmEa+10Z6nbb7j/4IzhwFDr4K1Iqa4j3I1v6MdhkpN51i/3F2Jtvj6hf+xjboy3XatLAukXL
U2wMBG8gMAbFs93eVatIrk/CA8j7+I6c6FU0DONp7h2yVV3T+nerK9Gq7lUmFNt/jci77luM2Rl3
M8aplu2J/kQVAvzRNTHzN2FMml0Cs9utr6Pe4XwCpNvqtztiHgQhymPMIWcwWgY2hZzFte7hQRxb
cp3htJH3L98+LXopNBuItNb+qW9kWjM93eLI50c6g7ziuuNIeYlbEU/vxG04uyixwk566MVqK8Mb
P8k4mVqAuhvvXFtXrf2AtRJNnBszC+SKDZw+R24GlA755qg6EDe0/kFwabvPOImc6lFc+44P+fkz
ql8zxsE2e+q+LWsU8uunVRNhYIo1Daye2Bwh1fHtX3kWcxHtHB75LHOwHy84CX24idCmC0bS96xW
qh0Wf+pn+G2HtGWy007tz7xsP+1AbLflo81Xe4bwf+9F49V8X/pvmd0Gb1FffJWSsgWNShsaFif/
see/a1oXeo8yCwEnVXDEjwydoBa2uDut8YL0EjN9Rg4KsVBIT0MNe9gIOhP0E+djQQ2X4aWX0G1Q
MbhnlPsfaa1jPE11RtArjOjnoWOsrsPYEk0TF6j7F+YQvoKadS6NfQfWEjb0LKaWJ05WsJ10dzw2
IYuezlr0gCgNf1AgqrooNFHfNWjZON17y0jnybYxFMb0fc5mxEEd7ccNUSqyvv2M0Qw97mnOydL/
FYNbeuFkqvcfWbaJjF92135gGoTmhrqEc6qHWPXGrGReQMQ+R+QYsxyErdcXoNsaI+eVU2QkZmya
vNtrc1rPwARm+R46YPJPcySe1W/1jTzw/Vr/3oZvdk9mDYWQy+K67/PJYq9AVECijwYIu3Dp6zlm
Y+1sJQn5Q7jzlq9fqjFrXbNXJjukXKiM7Lp3VzEiu8puPM1LCnNvkgfLxi4xK3iPB+cp2Abjyzkm
tqWPHqBAMTNAgl9aZRZ9ZAg4P1127uUsZ6MKywE1zKEPcSuSBZnRfZZWnt/H+2lua25/YR5kBDra
GMAOciVESyIxzjvrHu+VJWBQ4POowARNCmIBl9uDD5Z5BD3wzw8DYM89MkrQ1chsLt0ljebihmO+
nv9Gqn47WkFOZ5xbaQ6vhxhuCqFF5+oj0WrylKhZyiqO78zWWMkBcQhUFTG/0tUW5FMsPmrpTfim
Qpf4/elod1DMSqHq7WZlvOWtVSbCCLvII95P04897B9sqPO+p0rfjt3iX3yN2gO4LnrM/uxLUsZP
5A4u2AdE+O/moRaCdUAOAbcyW7LVY9qNO8ZZSAjSLJG37jsU3OW6gKnXRYfJw8dZDjLpZwsINd31
Gc+Ex8f55YQr9zYa1Z42mMSRTzSljKVbX5ZUh0M1IoolNorAckG/d7ijwIev6QnKy8XliyF2P71A
VeC2veIIoNGNjh5EWfa7RDV5xM5tZT/VJfPmELat3xLdtXhTp0BS5pFH5HLKF8A91xIYGgQY3aRU
sLEJhaTRccAYGFAtbEZrhFIQLa9bsf5BwpVGtsfdY2ahj63ejSL0yNzxKtv+MmawlzpeW0xA6zNF
F8USjp1IbyMeOuHbW1c5veaqS9A5nsTTYL1Fz6zVqsimjGL5yj93OCd4SN2FCY46h7sBOcxfTgWu
uixSu26Um3ciq5ApCL1aR/dF4AsNvTIiK4aUHe3VxNGtvKIqdcL2yfs4V3DlfgWXwXUeP3DkSHpV
/XRZQcE+CBnJ+rkhirE2JRIYTmRZq6kA/ekz/g39T9wAlNZB/UCsF/WlBDpFZOx1Th6hSAy7ZLbJ
6O3krp5m48Ax9+mqWAiqvDMMNCKDXvOwgOPAEYG6QTMRqk3L29lqMK9HuXmkK72GE8rQP6XVEFjJ
DsX5lELFaw5SYi5yQVtOR+ICEl061PTYUJvLHI8QE9kVbdypXPZG/+CqyL0L4H5yyXPbe6tJkp1k
63JfrdXVIizL51gBYAgPHjvsyilZWQ4Q+ZzomRijUCfrXwDD8csjFSqECrtTTqNaflbT5cgQqBp2
KRm0krWVgcnqtkdpcXQUFAqA8EU35+54l3oc+r2+UjkKsskduk2q1LvEOf7o51HWI1Ov4IZ/pfO7
T543611QCanqa/gKMfFAHM31DtQBPxyLfIGwpllWssoCnxKoVQ/G4iwskK/SOr4xyvuSXk8JVX50
UDmPgATLmsOFfKGcuwA3opnud1SteMA37+IgcJmn5WJg0NB11/Mum9KrDHbT3ihFLBVi+LSE8lSG
Bn45H+PhWgciW8U6DlGKIpAjguIg4vl/lLQOtDrjcYB0ozDVGYNp8LFMdgRoyvmFieQb/Kf01lMM
5Aa/jkRzNuMZXbhNdyrGw11eJ2Qm6Iz2xDlZN1qw1MPUDcNgy1Xn2TD3v1PLP+7HKeemW4SuZwY4
D1qq3v/VLd/Yd9BX7szMrhOv3BjIBPxZ4kHglhKiQuJD1VjuQIxCJ9E9tx01IK4PjrqH/f2sG3Ma
/SUottTB+HEifA7JY8cVukn8dA1oIOdteVDNjoyyZKG17SuUflmg4jUn7vv84LUf0JBPFYPPvF8y
Y5sXTAVHbQ7klYSWY9hlK4qiRX/VdXQlC1Gxowfqhr/jsAqisVnV4PI5bWsVpn3AhWn7ksJihKpE
nr340by38PADr6FbAtWgyPWDPjHJnS1rUmQVfGNQZLVR+Sk3DRQRvCiPnisVUD0SeoZOSlEi6mSp
wmQ+t+N09C3BdIyEFIntPTaoskpjAM0er2F/QO85GfaHIZEeA2ywlcnLw73PN2LAAsLEutt0S+/a
reBW6kHffSsyO/v9hoJWYl1nb6l485hbiez7OmavY2VMmbmE9PLy77upi8WE5HUgos5psizLAPHq
8lQMCYtmQBL2JUW8uxXHXkGUP9WGEbEGCnYyRNpQ0RWV7Llri+4USoXDGb54FgvnS2PQvNZDGnFl
anEbXmOfLnmWOoFyRi4o+BJeLHnFe1GxrHLV/BTeBFBrnk6elZqFb3ApYh3z+wMiC24lm16rQOPk
Uzm7D9zxR+0Ih1pQegXqnbgRv7hzx31PPZyoEr7ddSbUAnGoslARqv507FdjvH4R2KVw3WbvX0yr
U+G2EUh5b4+XznOXPUY5hmeI4M0+8uNECAHspYQOPP3GRZ6rOUwfViuiiI31OI2JgFYQv4bNfmca
ojYQxZ1H919ZbH7hiP3XdxoM8Jw5t2CcjMZ6NuygagXca2wCF8wTcEPcQQf38ok3c0zthQ7h4UoK
VJLvEPs4iaOZ198xJ8CqHFX0KF18sX6dCxaolwaBOu4twIDr9kWtSnhv13ZLR/4mwah/kd8np8tz
1BKqXnALmU1AEXCNNzCNHUq1m1tO9sdZ/9xgSDh3HPMwPvz/TYQF8WbQVDMz0DjB06nGAQBVHcot
gANEmt/jaS9kjPmwzptCk1NUyy5oKHp0wZ1lOrCnzKatNTY4idpAbKFhTrPfOmdng9ElFAixwo10
mgGtV+MRucWKJiyxThfsTZ8Ttsf462xDpMKlqWBHdtng1gbS9AUMNIrHGGFcN6skttz8uSDoZ4Bb
IBUjsu8CVwsWf0b9cUe10uFoFppBF09BHjI2nq6GVyPTokc05r/Dg3oB/coBZeNj3HNdM8PUNf31
7IiEU7pDGseiYSelWuGpx6wrDtpiuAilTsMNhragjiFI9Gsq0toyzNQ2I4+YjD3WQalyJWPD5Wy4
dxq8k38tRdufCPxtveXRegLfFu+9CSn3EXnoOCUJZV/kPDB2jPTCTOXVDpl+SyqJJAZKwxa2rVWV
LxTtGT1nCN6kms/tpWcsxerX6fWHB9RdjEU14hAcf6tMb3YBWZFvTxeAG2zGdMANneOnALvwZru3
S8k19q7OiRM8J92pnVl8Uq5Kfj0T8qxPBkKzPS7kd11S1NiomvQ71vsQES+ZPVpbzWrsSs/5gK1V
GddCGbh8KVWPdc33esFjSoPQg2C1uaXypONS3VWWWmzCXBbPLLYt0B0aJxxaeW7NbsKFegtxJuLH
hKOZpHhvvAP9D1SwCtel2x8H3zhDVyTpLarl6A/4rd2PrkFHxKdSNB+XKhgsu2/OU8ygt71HAuoV
1IX0nvdm3tsv20XDBITnVO8g228Q2gkKyJzqb+28gqYBwOLPNNQozwLU8e+LR19XOt/CAymEQ5YO
f8ZUS50vyhT4vX0/wW2CHTlbYs4U6O8yQ2h2C6RhzibckreZG+7mOJi/RInTC7CUKLOHaO+MFM8h
TfdUTXmaHFpPQeNNat7mkLTk10B1PbScea/Qm8f2bTiMgKmZXHMmwDQuRjHiFSIWESaw/w8aTBCV
1gRSM+kegrhR7uHuhA1VmfU6TTxTbOhj043w32t5+DL+jj4j9pPzP9HnP7YO0mQNurd8Rob9ASTI
flBqFYRNxrRH8/5v1S1EYPlmeou9S9NJFKoGlgTPDCpwbyQhGKNbg2cZbH7Pe/S0U3RVlzMSlrTc
UJYXeTeVx6hhkqIsFxjXzDQ+AF851tBfDqorLmxOX7YJJWcl8jTP5/hO5bqBU/T83MCTq0XCYAJx
acCIWOayLZ+zOqTNB30Id0ww1kNz+wC2fU2omCBqc9x0b2DdOB9//ewE9C3mvkqdVhWxN8KTH2Tz
j/3+bujBGCKPHp3XHg2QMY621H/U1d3Do471CvTE784/LtosindeI9G6Z6spGU0I6g6rimhGGiNa
wAkhjBPy9sfH74TNr7pCj1wb50dxhMqQwa8pFaitRD824h2gEFsWLK2mKpUh+rLzhqNcBRwozEv2
TZ6FC/5VgSPw34b//C+NZTX/6H5CBtJfgjyV2cDtZhtz94pmqhj0drKoiz8KqDp7y4AfYnLj49We
KxHzw2yaHk0uPrGlc/U3tM2szzY78VGeLBllICLQ/XJSag/aQUdSaaPcgpbTYi9MpDpsu7JT5s3r
c9OBXBaI3+4thQl37j6MsVzEjhNYUPSNRKabD8uLP3+PCWYQBsvCYIPpUPVAM2sZQPVrKGpP7lAl
ibXoNHafB3I3brfMrBqbiZijxP8zmlvAGnvTomZ39H8mzUtPjgJmOEDoYxzaBISvlL/3dbx27Mz5
wgAQtzIBUgspgqe2kizLhKOP/7NsZJFdRUnpSOZCysJw9Zf3zjy+tGCgtqHx7RyR3vgNXbSX6bkd
RLrKpjkP90V/bHTy4QtY/6jYGI3qLWdjJOcZgDypxRNX89cArvt0Q8IIMdloZ0/9fnEMkKMF33IC
mQb1iHTtJhQ8vxl+z2I4umKEAk7kEDLMZ5+g+beG/YkX3L2l3jBlL8OhCB5JXEJ5vrkJTfYEfOgp
fe96YWIEnqXgNTEqeVG+s0eBNB7D3BXZer6likk3H+nimWtURL3ZCshlz0VEUt9V6Y+l9efU4Fkm
xJDt6nB3TcoeoXnRKa16Y29BIHHtkrFR/nFCgtuYFeX1vCoMCupG495bJhLcAPWsUJmL0qgVZ2Os
UE0pKlkPJkUtG13HeY0wTPv7VrQTm6VJk56uDaw7BsJa9xM1G0rx4zLLUE3emP8YB5O7xJtq2zht
dccaj8F9eZibaHsVattzIar+OB8wYA7BuJfHd7MU0CuSXXYwsyEvxNOkvKCgpR11BQWEKyzJZgRO
wNxb+PNgs6JVzOAzuie8SH038J46Wd5KM1g4NwYMEXT3wrM9FOk+7HGeRcaXldUW4W52kznig9/7
+AtuZGggcTBAICQXQZNghyUYlqGEbJ8RSWGIpq/oSURw4N4pKic/h3YbMWJvWWyB9dACQAJBHCm1
ZaeH87MIrl9nfcoVpgkU4XlVuyDDMRkt0jH0A2xbBjGbGhjnbajqCXyvTYYJvauPcioIzC1fGVAj
zbYZSAgIs3m58g56ESnzboPatlv3q5zzCYyM+TkeV0DG+esP/A3ZgWnDldGcK39wNVky9hxRXyQb
P+Pe4fBmlavsRaF5yBkgUYPuMRYgkQk5ovIfyZYavzS4scDqY4KeEushemoSX92rqVIO/QslvmV3
6q1TfMHL6bFUpIt9iXQce26Fa9OvRHsRdNrEWDbTDaN2UXw8qiX140iqn+Fl34MzPO+W0JA7Z0X8
SyS7nqBIOuD1HTxAq1Y7TwQz3vdRoJP8ZbMR6wJBS+YLXgCpWlxL3SU0wW+5QluV2i0AlD3OFGT3
dJR/SOeHnIkMq5I1blFQVswCahYTIVfEvnKR2hezHz2Op8OM7yxr25L/ANQoWWRCmKUpikPiXaEp
K98K2+8tQ8dWQy3ilO+NK33aBiZFZiyYRHsffAYiHDA+1iIg4tSfwbBoxEREZIqHUXTxce1/Y2S+
4xAs7NoyGWwThV8Rvkwvs0UWeZzWFgtrNwYhB55v0aHb/gCh72pkl3hDQgNCbl8Hn6XayEe09LwU
Lkk7CBCQZxQWok5JBwU8F36hicKQJpW4pPJfzT9Rfg+vGsIKTGHAArOOPRNzWtqxAR2VUi4cdmpn
03hAx/ZhGCS5WXFPoIYSVyJckUpBaZ2VfK6LLOeQHID8zZ3nzGwm91R57B41hkJmqu1WRVi6xlZE
ZF2aIAPSCHfLPxbL6IIFDKDSwK0d0RSBHylhJI3JTDHVJ2MRUeIJZnYYQPr58xA37WCUA+8JJDBd
8G5vt0qQEYyqd88B5JXDQxp3Lm9i+5zn0z7UuUVDGmk+pKzxUrLZJzBVsq2U1EDUASYEgJmIKdBe
kEk3UDHqFqeeGLQbVT5pmhOyL8ar2KxUz+WBIL+WE2jphs7VVoWI67FPOEPKCfiYMaQARCsNY2Eb
iyxizP2A3La3GrcXtaNhtlgG+YBqJUFMsHLacfCIrKsBwwCXrzxxDSu6TM5PtJfcjGKBJ1tVKb3z
3FxRbj3EqmrpMEYlm4qWBAWhbtFH7VXHzMwCs1ygzqPkSRD9ESVcCscp1ii+W4iR/P8J4FhtTr3l
lLBmIp/QlGmommgHyiptqyt7nyzOnITn9rIzbBx1t0WqHssX+Rv4iirRkhiOayivMjqZfNhUUnTe
4PyxkDVQVZK+1n9WI7PuOhUf5IyYN4R4IFuWbuKOgS1ozGTz44GllKCVI/3lxcqSpLKd73Vj1d05
mRjV/VBir0ebYaDri5d3zQE34iAclAvP+BAyz3KTWfviip6geOb/IDyX7v2Gd5Mtj6R71t6tDUBe
dWEHS1JHR2JvHbL2wgH7V6rANG+35SNks2TNvPWwfCq8F+H/AMPsRF8AmpUiAtmDPf4mmaSuTXDk
ShJg82Kkx0bVqfw5o3sbRD9k8onUfP2CJ1oVdIkhNIN+2wqlGHdT0/i8SHRQH+CS+bCCEZBmFiTA
2OtijQgGD2N1Zp7DEjwm2B/IRLDtwRqkSOTd6cVpQaple9ARPoAMMBMJQfN/22dpRgRrNeHBTECK
UqQeGa4gDZwlRWyQcK6TS+w6zAiYJbyrwViyUxp5H9aNpruko+roYtDVtCzuL4qCGri7r+GVC9f9
CNwe+9wDs9gCNtwssORD8qfTWtD3OIkMA2J+GdUDc+l1j7KBvN80vSkkYg7z5ppkuTFVJpOxRG/0
UVpprGPZFDJ8GdVMZj6ZbIdo1s9a4wbQ7OjNoJ1J/UvrVvX4ePFLZTlMKWxIAsHImDfRA0KNvNu1
G+3BbHv5BDc+rTE+rAZKO4x6OJcDHmNKP2LcatUPX6l3krqomO6Z3JW5qgNPuTjGLw+VLpQmbp+0
XSYeuu+xs2OQZOZDXtHhQhbyzrLxdXJkwjuzU2tiBfNe5OPZhALCHRjGtj8StG7fIEZDzIvWhbkf
DnjbhDc1fDeafTWmEnuqfNdsshqrkv3Dgsz6sxlO0zDC/3HzoMF/LDi113wgPS/jr0uSVeiR2u7i
JdFkUFzVmuJ1HY6Nolt+EnrEjqP3/3XZ/KPjk449DyiNqy84BADzC12yNvodX+GGK6VtlZNWJDBb
uQ1/x3+AwBVcgkT24aPY8g13mW8h6wo5p1IBWKs2NpEptknmQv7cnbbBHBTpXWV/RoUdz+nhFBle
bUOL/bIExyY0FhlRA95OrVps6Y1jXm5o9tv9ovevOBObceKLWP9olrRI1ALF4yohF/P31MunREL3
4PYaxRXQRGvBnL056zYJlsNTzb7Q9dgsWjaOIbc+7j8Kpxbut/hWxGqQDhllPbRu6L+V/OZEawkG
hcL5O2OSbk7RSZWDhJsxzGyLTwFZIEhOzSaeMZyCOeQFRrFtUCycYs9rlVgaRMHp4n7fcmxbMgxJ
Lt+BbEan3oGSgVr5AwVsRqyFDkC6HXVNgM3shKHYGAMMeiEDsOMreVZ/xaQKwW61uVc4ZVWiGXci
Lg8/PwsZYz3GaFm8oe66+/vYN8fwLRrTuVMFBgxjK589iDL8hV27h3M8QxNC4sEFesLOzRy8NIhL
gPY/fJu2c+fW+m5CxU8AepgFNNYjgKYD1vAhFlMCvMkTbYXYKdelmsZnGOBnOZNypu264FhMiX6D
97/XNgEAemmN1ttZPBLMq1FjGizYXgw0J2oVQDqWK21pQjl8ZDrDJwqdCJvI4CkSpHCIwIOfalut
VJEctPACwcyxagna73+jUHCGurvtUVC6zXevtNCH5yxaJc9JMRHikCDSCDDrlI7lFbfCQ0o01amc
36CPXDVqKRVyRhxvr2+REtldH+OnV8QydfGP709dZ2h+1mlO9Ks1ge46upU+CgcwUeXG3+lpbZ77
tGJdEOF3T6WUqiIDv9MIUlouugTbX1J1GO3l5GswhcPkxRokysfSufctwOq2s6GZYEnCD60hsE7r
7pUsP2Ksi58QGfN99OIAkPlsCNjpCN4VC/KicuvMvJ5SD9xX6ozYmplrnvgn05pJcwO8HrjHA80p
xVjuEarbSOS1NnR9QgwwnatYYg87tlOzDgqtqwVJg4sKUJVW48pwMqQVVLy1DPxMhPrMUq+uZu8+
3FHLxzAa09OEpwfTXb0INb2LEadY+wVG/FtTOVTgtJG2HB+6QBCugvIFibWAF1plD3KzT2dXGVtG
/QiUVTlXXp8fKOWnO0Be3W+CPrEFibSHb3ve7vxLjQq3pN0VLr5/1q1vZMBEYlcq+A0rlseZRS0q
g0I9WwzFLnY7YEo+GqDq5NTilFvZgLBBmWwD7fH0hOhs+E1zdN2N2MZ8dJlDVd6XwWcsrM5NeXLS
VIocM/j4vo7T3o1oEV1bwIY7dY/sURk+2mNohzNj9yrfWPqMz/7XQaD07JZhsQMm6puw1MwCg+nI
JS/paevQeQwmPMbArqoOOhJuRlWXZrLrBTpXsZcybWn7FAtLgWIY/xEb7Ig07gHzsUD0e1oGHhRy
x3cXqgnu3NkAcyYl2gOFY4I91e6sNrx5damOU4GnqWdQuPh3GCIPbAgw4fET8pbFNuY85jSE6W4Y
3Xeuq3/RrmwEhK/IFv5NqcMVX+BBqmD8YiBdnmzmZ23TCov1xlz88r55Zs9TgZPQbNa2QS7AnQIL
R6s9hEJMTCfKc7ocGc189ADz6hdLL81BOQ/ex6/wCdB0mcFAQpfWkx0WZO4ZbS8YGX8Rl/7ZESnd
NJlLh6bbSnNhW/snrVxqxn9fHPQRJawFgmuuSH/FEFyvs8qMlzn4+NYUqh23MmksoGP9rxCcpDZe
qqAB/yl4jnktF+4ui/PnAIPBhmAVcb1hCZmtg94ttASAyIVU5Qa2KOjlAcBa6kyX9cpclmHHa5Nu
KYSab6GPmF10WJ4k26vthWNsxOe0VmhequpEOI3vrYcrdvrN6YtSDsyI9A+RWaq5cBClRfxoS2pJ
y/oKSt9p+8aV1RUnyAGqMMACZNMkeA2ooXp2LBn3LaTGakDtdeUgFBTJSVgr2ugz0tXIpho24ZQH
S3dNpXaNV5UHkvuZz7cij1C/N5ZdY4Owhgj+57nw9RmLuWlQwCZKXR0XvzBdDCyhjhroiRqSafsX
Hn9A08vg6fejLY1cBev9kOrqpgZVq2k6gS5Q4wMkjg/PXzBK68L2sK5Dhlgm2vqvqNdMaj32BNgO
k+ZVsxge/x9LpV01r2VpI6lz8hqixMGnNipZdfKwQ7x9HAHCuBjb5jevnShP82yMZwGSmij9tBNo
gs+rcn70+os/vIQWQVFQ74Wv06df4hxd554UkAx/O3yOkTQRRFBTlOsCpP89gVooFuJWUwg4G/KZ
lZm3Ws5J0kx3jWZjVlKqCnS20YTeDwEBigR8+04tMzIx/eP1sFJbY7eRmbrKPPssFskDqvDI7MT6
/JAJoQXQGuSIL1pvHp0fJZR/mfo0gkHKE/HX1pHhYhfT6qSZ4pQVD/ugm7XlUkhkvG4xmHLQzFm1
m+ihizWQP0oof1XR8IU1wormfRhZRRbMVnL0AP2qvNCzX90K841exRsCjGitH7iHC7hXmrAtJI0U
gEa5AQ/ymc2GTz10BJ3PBkM/9StnJe6EOrGWCLFhSfIab4/8Fjh11a3mjAmj3KXwcR05DtNNB40P
XGGhSM/eNSYUQQb8y3N4cEsAbZezHiopHIqehBznhj80pNLS7w7xw2ZwIVHrDJKbc4aX0QvUFwCU
1aaOJqBoQlq9tqcRpfBXUpwLj0nRLzjyzpYLmrmbPf/bWySifRzC8VoUaZdZ5ACOkrcd9FAOhkiR
pvlqRKinXQqFfaV4QIamAxDEm1SwzlXkU7HeHehAyu5T5dmEi+r6X6vGuI0A/CqS6X9GMZ1HiClZ
aQgUTHZMlvcI/tI19u9o9hxQCXjSQ4XVoPIvQauOfVFSAn9WVjbZzOuZsLsIMyNgO6LaMcihsTqb
zdNbVCgexv+NFBQ/RNZe7xW7/VmzVccGs1a/Xq5e7kWOkFcfc88wyVgo1d42UkEZyC4VzutOTrU/
WlUellf47qNqq5De2+RMYKp7oYUK1Fb0lnb1lXa4YGw2hBQcSMdEEQHShHKD9FstbVS8X6+L6Co3
ZCJ/a8nMEeNxoqxYW9+q5RBi4tiXdjwZ2VW9wZFr70dhe+MzrZxvBZ37W+/qXo8+yuBCOWoIJQp2
TPg5tMOAYOYIy9su7CLzzVaEI9rjHqHHJn8y6XV4PZZaHDI1ikfe+P6kk74oI4RTt7xlb4pNflqs
t0lQD0EfPg40kX+f/d9pJfruZ8XxrBbb03cBVE4r7gT2mjp/hryFII6rw1HM9dcArvF1D2Q6eain
fcHcsNf1z0pa7RYlrCM++795kuJflTl4ZIFaFt6J1Fi/JRjnxL3XsKvClBdFqw4UPB1Q7omY+VAk
V0W2yQo2OAwN/Gkd3H2UqwwWkToUbnwbrEj/01lRHKd2xJcUIU6TOdXAJsFL3V2lcjiM8oOGokJj
o47j11rxRbG2hgmMEp3KAMzV7OK4ZqEk9c+7bbf7K+ZYDaeywQfIWHIr7rSX4jRCkRFYiGA1nNSY
iirwF3SzQ74nFRvt0wlRh813C+ZnIJDzo+YOcDUBJy/YliPUWOPbtzEElIPQrgYSG6qPAWI3T4Yk
TXnBKcD8o0T8vmoBBMi/qc++YcKgD4o8MFG7LsCT/kB1I6irTsXOlqdU/Bf3BaGc4xZ/DVDkQy74
J9g0tFj8a2SthlitD1DU7CM6H5P7OLCqn3n7jCXnobNjHAOI/r2dt3Y6mAlrJioRlcqYTMDUXlzW
HjKwYAVxVg8fllodX2M2E61Uwgs1snNjtvidtcQvqDMUEr7n6Wg1NsYiurJntIIyANc6jdZmR4lk
dupQ5LwJevrQ9EjURgAoM/zY7KrKiDayZDgugoTAa/P9V9AeLzOnImk8KgRR+pURtDvfVNhBXvYO
ObcAqIG5mI3xR9uS9HR6ELwLd8RapxmyMNV6xp7mUWod6Yo6rPMRPGL5FZQr7AErDDWXBAmmOJpk
R+/b6QP6ke5wjB/pKqjuk9YGfulb0+uNkbTHNZ417nRfxNBqvSxTAmxDkIux7X2bFzvQWnuHO6Yj
nKXhHmW1Bi5Mtd6ne9/vXP+NqtAGkBFdFOJLeNUi7ZW0cnB9JHfLIo3jmUlvkIUJ2mbsAj9FqC5/
ysHYxvQrIUyCY6UG5mGkLlXbbZXE2SLzBTQZCWWbMqlzj4TwBp1drpYep9dNVIkrN/f2VcUji9Cu
fYwW2/2oLIXXFrR58RBvAit4ZlyiudQd5iYRzj3e9NHpu6FwjJ1/uYPwcnsPohhfQLvl7y1F5mOY
9V24PY+nrFXmmgZv4D1npnQJn7P+PoPaOEQ/0wFKVO97YqshC9VWX78lY2sFCS4ztw9lbfn8drl6
wWTDbnPK/62v0Lcrsn9rNfP4iuSor/UxzIVEEazjdPf4l90wwDDRxYpr29Jzv21Qwoidq08IXNU8
9OJrMOgQl4rU0ruEqdP0ERZ5uic+WZ+bLv0GGJIyOfj8D9XMpDz+8xtM9PbV+mWtBfK0WIYCNNiH
MXBz9kMtu0hxmA0FJdszInZfaaNm8Mco8xfTnGE/F8Gok0C25nKyX4PSLGrzCCYpLdZ4LLsrRW1e
9I0d+duA6DYzJKJk6wdCjX97+BIH/0lJiTu0xqekh8/eR+jIBwfq+Z7vTZvRY5ONqPOHy0ZH8UaK
cpypWC7gUOVe+6/SqqfdzajVCwg55DoxnwhtcmKHPiB+Vrjjt80id5FUxZkTGffmFUQzAmg/CWeR
JyrxyUaz6oC6H9SUJc2bnXEQtyH6J7yC5WSHv2vUokLVV4tQMVvqWxCw2qAb2jvz6N5HyZ6HUc0l
wxNUUeM/HzCSpLZ5pJzec7eg9p85nKMMlS7Te6rbuV5hXFnusclR+wW4rnLtB1IzK+Z4tB6PO1nQ
ZJWiGx+yXQhjtkRElbYlZvKlbnJ9rqYtgtufTLeTzlNLhy0lO1nSir/qlj7r/vnEknWO0NPL09/a
xC8QnYx4kpbpnca1nwt/iWYSTca01/tOquMbDdUtf4eynBxqEJ9pvb5JdFgy9PZqE7nfniUgWdeO
qTFWT+zvTGf2HSt4GMGwbiiylxP63RwhJf5HVTg7pKluo9/EAH84lgeThO2bBYo7JuAQAkxtZ9YH
XWt5rbp87Ormh7iusmuehFc5BXBmkYvV7kgpFRG5/fKTkcSj1IzkuCHgudtwYttkOpuOnbWMV41c
YdcYUJ6kZyhCCUH6gEwqnKBaNyrcds3mTE6bEb1efyj4Pq8JfA1tnPqRTZDmGluOOjUapN/WAkMg
caeHwYHqWTDNeKlk+QNZ1dhQAl+Zj9+ukcAq7/hWY+C5iwslKDAWjEyEtSGXTUncwvSDce1IVdin
8xBcVU0/pmODcaSQxUF9iorpFeUcqPqnJ1sCyDOQrxJbbNpNq1xgrf1NYHEJm+bl5jHB4aeE/Urd
zeAOUMaVoa852qDfvH7ECkoLA/MNhP3Huns1GgItHSvU1xdE1UIOTg/KK7isIVrXgGfZQDfJCk52
+HUNTVbu9T3qAlNj4nb0+XBmIm86ie4qBa7v9sSlhdky6FRpRiAvXCoJ46OIysKKd2WVOiEcNGjf
Q8IW6A4jtIVR8x2dK2ad9iYXRLmTBdWsn1QnCDCgmbhguGjm9qPlhYxTQKYDJXshKKLcyzsO1Oqq
RTs7B3qG9rksYS4l8G8baXZv9mdcHIgP3TSm2Z4BirwgCuaVh5SlM0SxIv8M6byAwlQpaF4xsdV2
zFUdoDqTmyI2uW+tK0rqqIlNjbad9jd+rUIXI4hJG0WNANyFNkhuCDo1aJShozSa4X5omaOphgQn
czsy9Rt9dzryBgIEXxtP+RlIz3niFO9RqktzMLMJc4Q5l5TaQ+PWvVNAn58QDpGo46mVZQCDt7x7
W114UaX8kkQoXDNvZLbWY+i2utKmJVJY7DcMHKxtC/Qjb1abPsrK4TGhcSSJZb//dLRss/pg9ATS
gxUgl2kXfV0qUmuUW57gC/dufYDCPz9oCDoiDEeCQtyKxETQx+mKikFSkAYKZr7IQJctsQhg9toV
RzVX5AnofcE+Rn6WIsCFN7+gGiAMgobMwZgxRxschGeFKrIBAXKUpEc5Lfg+mCpFT1wdpdnRXyyQ
R5+lSficW23bJw8mTRTOwZDSMMijEmOGKmljmP2SAhSu3FZdXV28x1P5BDtqLb8855dBCeTyC3kL
G40JgMrEfvX/Ar0AayNSBu1IDCLy6LjseSoNWveq9I7CwlsrGEHL+fCLH9FeV86KDsFoELGvR+69
umN7aMTqi/l5eheIiO2i3ZOSVUjDlnwPkQNNZxwS8QrW39ziy+ghAJZERch0ucWjKfZMINNmw68f
HPz6iF1/HQnzajaZYyrW1aMz7QNf5jYKn3tQSJsjaeY1OekTC3RVRSvt7qnEG+OIM8sRB9Uw6ePc
5VXo6Lu3kD9DnogaWzbYHwXeFkKk2ZRmTXTGvT0o90hG2XgEHUNBpd0OnMgkAYH6QnC4MMFJegtz
7S73W2i9v8JMdj0mUdck/6YSVAm4vvaHx8MCOonnxvBGz4spHjjY1copc9LTF3nF30rvl6FhjMRU
5b3PnxrcFhU3mKskXehSuIPtYOLsR/cjqFq9oogsFhQwfyMikL9ImWFbErtIiQf5JIBxe0f32Jnw
dKTiM4pWPIMCcEY8qbo/vQg5xyXj6F5ADlx8n5Sgln+7KoxZ+t34uuHckFUkfJDeuxjOEq1HZbQd
Vu7jlLJesVN//WShsuVMzMhtCiZnr6d7GTgs8Y/5vH1xj7lZJxJP+4U79vUjZi9a2bOq1i+iOBpu
LgUju9PdsFleM93JmxRsosyH+lyNuC82MJ50Y0eJnHURY//iyK+LJeNGuC+nkyc/PM9pjcQD2KOe
sf8TzDRHzhOw8kzOXsSoGZfTaBG/4SC+GuZ5i0C2pvjTsFxLI24/xYBjBnheryWFsQC0M4/Z88zb
z2v/gtLeb7q1/l0ELVMmBsG+oGmNyuDv4ZdvzFTHoCEZWkD6K/+c8XOyMrhBE6lcmBejc/I2ZRAi
RtWxgNDykyu29UoCFL0jYTcl8OBzw+R6wh25a9BAYZnWK/+Lb1Q18ufoIEFMumK9CtgujtECspL/
k1ChK2U81Qp5Y9CEHD+u8Zli55nmfMS0WhIP+0US/x6/c8UCfY45FJwUUI3lsqwUIYf0NhjHqbu8
crYtfmb938AymH2wRwKxJbabIlc3GyQtBOdk/AYbt57Lh7+q0/pEbgpU4LWaSp+Nwo3n5E3RMnFT
Tk+92Y8tZUsGUCLzusx44okHE/dUVkJNAm1ppMLcXb0i2ZWGg73ZsMnNWFGkixnhnYX0Gs8xqpxa
JNrx/k4QjxAOqhFj51sfxKYzYdO7u8tCGnYo6eH/Dap401pTxVhuBNvGFo20WQLqMaCtOQ/lHCS/
+rz6WhybpicpSr8g8le+bInT606PZ+VCkBsyUJp+7ucIgMwpGrJ8RVJj9A0dYDRtafJS/+QRIy9p
1D+WP9NDvwEsBSFeGtK5ANNW/YqZZ/O3t9k1O+dM9QhIvEKDxc4tHMib5Boypjv8xY6x4G8s5IPp
bw8F0zlZXCetwysR+oi/P2JqdlByydMmIRJGxdNf2TW1QChQy/29m6KZvld/NRCv49LwhGMg7O0F
I+SNUikGd16RGvn0dr5wM4KZG5g7c/SLZ7v9LkGbNXi1hZTrpFQLmNUpkVnEJxSej8lHjJ0WsCG8
Un11tg4rElzNIr6jj8xSePrAS1wMs8PASZ5FsWz1xt6GW7bpKY+doCqA0H+9N0/YDpgDUX/4T+lD
eHg0NDg7CQatqSsLU32rtcTxdqv4lT7b/RKJv+TFgwVauOgWiKxILy01qJsl4RHnweYvbe3Bztsk
UhyFm82u+YJC1vKsIT3jXPh+t9J73aMMXpBJE82SSQc4towm40K1CpdSxIm5+hlNv4pkJ+EhBUQb
CG8Dx69YZgiT17mGY/ttyx50xXsc2NzN+n4QXwB6ZdzX/B/Zwjg7EI3D2xFzx8Ma3acIo1AGI+Vd
zIW51xX3Q8kqfvgXWoUPen2dc+vHiLH6u8E5knJX5ey0vMF2QVeqmLu063zoB3G3jVNQtJTh7YO1
QjGr6FDzXyEVN91wWNpJkzz9pCZLPoeEY1pfMVNU/kYQVGmd7TbVcAuf6xVTJvT79BalIXBpTD50
Dnn44Gsc2GRt192AIUpCHQGZ5AGWgeYCUTHyjiFm0ep6Fw8d6JSmrshGConWDA4DdhfK3KXF0UDp
DMt2zD09yJAT4wVv7Rmqrv86CwytNdT9ImYJlkT9yBPxGu/1J99D3YSLV087scHfuXv6EoCG2gVt
AjDgy7pG48N1Pox4mMOx2rz62MH7EOJdWRJg2sXSL69A894Drkf6LzanWrWj5xY8mJzkOH1Fg9Ad
i17Y2hOLA2wJbNCEixEL8HrI8ddP6BcUkx1b20y7ZL3SdYeKqKnm0jR8TNgsJhZjSK6uZPLnAJsc
7wXmXVp/Q+6vEKotw+AwwDeKCkXb7ALN9NwSf1wqzBT48YTwoa95I617eRZXWdLNDIMJ8MzviVnq
bFihD1RfoO01/569cAX87FSTNnX5JOhBbmzEKy30hZ+25/g290vZyYPgMVb3guSEZK24ib/e8cpF
+27loSpHe7hHfYi5lFT3804WGYOdar46k/mdikwB8XE59ENDTx8YHoZtAytcfGg+zAN2wpw5JTsk
xiQPzNv00UL8jPoN/X1zLIVWJCwdtHKcuehjwuRY9X798LugKu9Fv8UOBCkCZWa66fIPltPAr/mx
dxvye0MFNh0K2cNonnxEVRlEsc68MBuB5kkv+9jA+6nu+byHtzv2++UluiCYsyi11k0vwmsL47vD
iItTs3jopVDWYrue9T5epWXyg1pQg1LlrXJN8oiXXDQUdfmknrSaeppHjBIcHm7rYGAnXLsGWgLm
xqvharMWR3jB9WXMv1EQbKdgHiPFhEkXvNt89VPUKLBwDuJU+cIWAVambGHliqQboetbRMTLRpMO
04FxZvZiZ3SwPlnSGtB9bfMc3C+UajUvpFrknXCZVJV8nHgWUjfd2XMRTpm/S5bXJfqQ3SruMNY8
xRK6lAyetJ7Qn6G6ydcy2z+Pp8BLPI8j7qf1F1JJoldc+acHoWq6ciZ8nl6DmMi0O+XQ8mxJMlIK
ql6j4TkSgWjQXALzZerNmxCsEPOu3s5nO9GQ1SAT8unQvvEHolHsYc+IkiWEfQCIuZlKFUQU6Qu8
IuLL05U56yqrQEEwF/ymvz8UkVwQC4Einkt15o5Ps8sE4Bkp4lYbuq5UKoKHeN1sA7h9H0d/lWV5
ZH/IXV8T0i7HODnJo8Lb4odmNm8XT/cJmlhFIQsb8FMqDzGERhwFdT0PncY5EUyH40VFvPcpMK5u
wqtaY7tUaZL49JrHatMYDj0oNHl8ZHSas2XMIYR/a1I1YyhrGNZ8raPj6YBb6v78yU/zv49Ocw0b
ylMy3axGlvgUP2Rbq0tJV4ECtTM0vWBmZkEwjdszQXm8pWaww9wlF0tLouFzEQX0fAdBRVnf4wwh
NX6lu7q/cHF7PGu0NEWcGv8MwVU3prXR8W9DNUNIK2LX8sK11/Dqbud3AO88oSoJPXgNStvFDdFt
LW+zFXu0OZHJaIhuNYE+7QovFQq+rZB/bSW44nPnCIlqD3fGnM+coBpNh9OrO4/JMmVugQ0eqtAg
cWk48XK+tVhx9pCz48MwXxiQ7vt79HpdkESjnQiQeFiHXP6F2klUbUaVfrm8Q4jOSDw08uGaZkkV
906BRjuHL2O/Qz+6286j+DAmHG4b02PJC0YL3R4ydcEhdbUEtsG7680N2fSDCjrcpUKV+I5U2cxT
WbYTrmpIPBf4oNHU/CG3rPkZX7U8u+CZh1v1B0v54Tr5ovk6ZnL3qFKYqMhdQ8yArsTdPRr/VkJt
QHv9Xqbx5z9ZlkKuBr9FvcVJ8ImNoBrZBLO90UBs4FCGDuuS065de4i71H/xZR0rOH1nYsaQwOvm
GNVzUWHDdUuKI7DhybRTaC6/NmJrDBP0aPL4HHiPwGXYen5xt5XHD/Vkz+FFDaGYd62HTnuHR+gz
oB7ktuzMFWdXN1qwY631azy8YvdTQVvnQj2XM3KDvc6wWqBUq/T6vDQha2rObhrdbOpWaKTAv/lM
n3D2qV8zdw7TVpj0rX/gMj7wIvF8Yf66MQ3iImdNTM5HepOM0o9Ft9jIxmcUxjlMO6sw0fqz9nli
Hy7R//6/wtvptx9UxKlko9FgasOqRj79sKJBGBVGei/Mz1RQypQXjMrniE+hgye393M1PCkA5YMa
2R14zW/7XwMKhmZqvJqmirln1rWJ8BNG5CnCXs28VcZy4pN/ccYWb7edceg1MAzU9G/lij2CbYyN
2mDdpoGBQeIaQAWmbwAjrhmPglNeL3UaeP0ucKv/1XyjTULbxUmkx8j7eSJk42JAB7CnCvKVRprm
jAzMSSEE3XV0KhkPlmGcdBWjuWbessdPVhBCYfwdx6Ybfj55MNI6XaNGfnLSOWtDSWkMlas3KfWw
cFpccn9RXp9BzreCaotMQKqZcuOkradsVP7qFfHi9YdfsYlRi+rFf/ia0Hr9wHSt9ly3l2M7U6yD
uB2z67Y0ekVsU0P2zY8q/PEPuCtXNamAJ4++is4yCD5p4O1wZyhdOBDaqN1fAHSENN4hJbV1JJGZ
SDYGn//bEhiHS2pfAyHMlXVhzR12KN0udK0nve2m7KP/h1xGQM9oFhQK6bwH6K1KCMxQKmZ4os6U
ZqyMzxWalVKIg/k1hHyiUmzCSrMeEflO9FCx3nGCiI0FEO3YjyFmgk/wdHaEDs8851IaX9cfRyTg
oj41HyDZ+uwJ9lnVstTMnI96aS/aoJvXDRSiyJxH8Lf9csZakJUQKpY9mVgOMRjPS470mbUlDnma
eJukTqn1NHi+JHx97LFR48e8AmOZEvV4Z4HD+lQJRYQZbGKdGmc4BTTxRpnVXF6IPuO58wrTb9e1
kPcTtI0Gav9e1DRBL6V3zC5bU9tEXg4gPdNuPWnE/R3Xgixvabdq597vbhgOWcNlanwHewUO7x0M
Bf33mY9UNxdYZ9BnZ5YFhvk5up17IYjmzZBGAZxKw6m4qlz40D7j5zT0dfyzszKLUAFlC5GEXzVq
iYgZyNZTabpcZD53byI+HHD+x6X7xsoaMcH77vlDgtVMy3P251W+ZCLVy3gjqfMwBiVl9WM7uqIz
QlsIjkndb2QP6g/0Jj2TnVfGEv6EKFba+iXBBPqjYpDcIPI7orrza8WuWbqJFF7sA7ZVBo+fKbI4
5Oox5UF0+mf7zhkPYjiwT9t/zVX3DDa0XouxDQc6MbVCLWfBurQGe9ib/TH2RgCWs3Si3mPM5cxO
Iom2S6O1ulkmMqmcjyDlh5scp9Hz52Gk7FerBBWRpxZz8pDnu9RIHVN0e39XU3FoDomQWQ4LeAb+
9twunL4ioiTQP/n4aHK9S+P5VNwVOVC2gcGornVQPX4k3LY5tx8FEnFpzgP/FQrylGQpKPzxRfqE
tBw2Zl8QckvOvr83gr2D4Eu/Ayg/wbc+rNrA9J7ArlAtPgrFkqzLS/w7taAW8Qc0JJkyVUsgmou3
AgzMJYQKXoA99GH09hRRLk51n44DRkH9FPmoKMvR5qMxzsl9zl2nMO4n2IqUTDwkkU5wnhlMf61u
Bt9EVKuqVABbqPtWMkyxWRQ/xYY2FZmUKms9XmKEfWluZlNC5VkNXl/H/ZJ3oYnfN7ORCbrKPsTw
HwESTxzc2XB9Kkc5IFKQkUF7htf/0V/WZVJiiOxT2RqFQvi8S4w6mMfGng70hRx65szBYV2xIESo
LhbDxxA7vSIxfwnCS+pTW3N+SttFk5KBpXV5/EsQ1Bwkz3JwPRA+1zan5+Hq/hAONPmS8Z4T2kp8
UK1QmvDyG+d6Egdfpp9Ltnbh3+nCDFfF25DXkUIOD9UafV9vszxsA9ajJre1tRhSHOuxgUdua0I+
rT2cGzD1sFl4vBsPUNnvVLuA3kudaatIQDa15GqNntogOVx9Huau+41epuB2nb7mGvmyZUdg9oKB
Gu3r+EAMzGAM2tlK5R7Xm2DyCUFHiVUL7LDKR7nuqCQzjnsAhQHVBde+66cisMXpLZPWMiEnbdSg
wyO1zZclqeRFU05VUAjKwC7p7i1ho7GfE6liQgbsYQacLXYoaJNuDHBUlQFg7SA0VhpOjutDzdmE
cJmr1X9bzdvwV3icYtHoqINOkeyqJSk5i8xHyqCWvn1t1taGmR2JjftuM+IyhfqWSPIEq2DiQdvz
+YBGS4cYfP95/aUBJBhwA3wTxs/9MCus6c73icPj0knp7fyfzlj1D4pNs6wMTjCHsYylvkr0W0Kx
FCIq8Fa/R5PhBodju9HOkUD+9PKiKrBzQ0I1uo/2quXvpe/jtvphfkNqUPkwxa0zPNh+oAWkLTRz
OB3uXvxhCvO3r9Hvmv/DZjhK8/3JQ8W7Pe4GoVYLpiZPWsmqPThO4OKhTbDUdS4Pej1I6fWUMDQ8
USelv7RU22WSC0hxN2B4+XeFtPMahc6bkJuQ82BwbTQ1l/ibE3D0rJQKb1UcFcX0mpTTSfTXnUa0
BA75EV1jSEjrOKDfS9yrzd0XxLUg24xaCYmd/4UGpdiFXi4d6W5zU90CQpzm4SpDjhEUx5vkrbVA
3PdgX8IF//GhA7o8f67bub3yOfQ7ChwIZhyuc8HVzuC/nTkTPcLTQcsNrk4sxbvkLmOncwqAkZ76
gRKM/b+cdxkLzZY2tEs3lXEgwHhJ0QOlKNyVVCdJMVEl9Ta2XH9KpA6N0nd9jieNbAXUoG+gGr9c
tyBhYkfeFy00VC5hXPZlUIx5blmYZWC2SSw0sD7ubYeod2b/kpZXIo+7nZa04wn08xG2X09tf61y
rOKlrL+x2HR7BEMwHjccgsyb6HNp3cPaAei1+OKwAFdq9FN8qbpVd04AUm72DZ7QWjDqsSSCPwYM
ENFnB3X9vPDysPrZvX9K9Rs8LfVUM87DEGUf+8cJr8prlZAc2b2/Ea1Vqvk2vAhQXvf7TBJYilCh
9QuVpLRa1wfGdZMBnMax5MzCHnHXu6aw6ohgUjm4/alwEGcSXUWF2XeuprbbcAB7cdjPunUAineE
y+L7T73BNMpU2mA7NQRpAhwM2x3erwhU17onS9nz4uCrwO037WnMYHNBQu+V+0FVo5+JgM7BV0QZ
pMHqKXThyEdSUavMZxGlHA2kjGJOM+NYspX4tjRvXaza4JxSCkAWdfFEE59SxVsnjcPR94yGsyvb
RFlNCkLCH/++UbwHdZkr/ASS+IX7fo33IYPX+ogejFbUeNOV7M0+VdS9cs186WKpVRGVKERGUvXw
xpVsgVa8mvhQHkCFc49xH60SKQ5c2OtiO+L3zotXkOGIDGo05bEIXJnHoa3xSYJcPmO5GkB6UGBD
HIhdGRk25ekDBjRnVqeRZIPAPjWXqF7IBYcRrC/OGZ1w3peoSQ3QG9Fo3yLyjo4VCNzP4fpAf8iV
5WtwN0qT7NBzNSXuoSM18OvBudroHWzi6cp7qttwZhGMcOzAUDrvRNVm4/u2ZMcbGVgRhU/Q2bEN
GiKzQyBQE/E2g15r/zepQRfHqx+OOen6Co3wY3AScKbmH7xlZtjM4gK+zkIPcSdH9xiAmceRazay
NA/498BK4psyjJLGR7zNf6hgkYPwVAroJdFFEdST3Ht3aF1MFSEtp6IURGlfFWT7U3S/cyM/flqY
FHeHBK1v9IoNYzGFXV/bVAA+pTWsGy7wME0TLD7sWJflPPdNV9Hti9Q5IUU+xJ8eJz+hXYabg81N
ZB3SNo2soBAvzNRwc8X6wsgHr3wC29MDw2pHKUchoo76XosfGVT26xGTirr3LWZwSNpHbYcDlGm9
KAi/GbrXkE/XU00Qs6q6Idyp9pRxI/y+6ArQnKiFZMyWiAiHRrGXxVrP66WDT/R7vMHTO/KeHP4w
tlXcmRB7RclDww464iKw3W/rR4DBVKaqa9CBFJyyxrwcXrlsWDNbu/ZeJSxQgGHYhKpggC2aAR8q
3gmlCmI1wVoTyUy+CYTnKfuzcObdg+NiEvjhYeoI/Bjgo9dub1st82m1FoCGaKLr2EMk8MzU1yk0
bNUjitIl/HgxCCDxCYQ9VVsLsrYClgMHO5gLVOlV46ahz9+NIZIWmPAWXM5Ai79bCGX/ry9wf7lW
S7VkwhiOjXUnW9FOAABCnSLPz45z3c67D3m3w2XoPyYr1q2Xa1BZbfVYKIt4PQIGBvFPcirYfbYX
zqpDcqGx8W8xqqxcoZU0fM7UX31XaparP1Z4oC09jJ36WMHGvnBI+SQmBrGJT+18WPK8RQ7h7OZA
0ZZ1aGXquAuatVuR0CNT6B7N8sAs9LR7MfQmhJWp5ZFvIaSDTkg4MZLBE49/DxuNbJbFt82ysB9z
QX+QFp6//BX9iEz/MCw/JFxpLVb0Q3rxmTQcF1UkRdiydJ8YKZ6Ddkk+LiFGuVuvfcIS0nK5fIw+
ySftgsXs+kZIhTwC5wwtvuVBTbeYE6WCGHJ/S0shsOoaT/JhT76BqopvYDYAxgE6bewV+50bs9Tb
4h7QCMGaO2MRMLgxsbxkmz4d2AmzLGd/+6FCxx2N2IhpDq/fQFwCy1nwRs1+0CdOmgsrO/S/paJK
oe1mBsAviHvCEk7yYbVMjuQ2VNbTqKuxtqjLEAdjj2EphFkehLByvdAAILXy42NRwRg5q5uhAxdk
G0Yqhrugatc7Lfjti1JAU4SZqp+BbUga/oFTwRGLzRLvucDCjSHmrJsRwgt0S5r3m2hDYzadNGry
WQsyHjYBG7KtTpecnWpEWrNKH8xi9V3OL5jw7Zny3bB9I+UOsYKCjTFrXCox2uYpH/CVasVDWzQg
JEpgTWcApLeYeyvbrm+n/EQwLC4GmTABK24DWo7Mie9DUhnhFsckCfWr5f0NYJDeK8SBUXwJdPvq
yxpdr+iuL78BeWvicVGHq6TMzShZiSLMqgqwAjk0t5vJOoYhnJ0WEL7LzI1CXoMw43dKVZr26CWj
uxRgwMjtTPmShUtYAW+m2C0qaHk2LDt9Ix7DY+HJq0qMANEFVWPeXpT5PLgNRV8fBS2Mv45okPvG
joCUrBT+HpYqiUAm2YVBzBw0TwBVm18lv/wqe2DRAXDIMDzGZt7oFYIUVqY1ztAhyu+ZsbYpevFH
xyoBXo+fMzeNIyMblM08Wh0uQx7qsHTLX0ipQDb9l24iiK8T5ZqwHlXcjhVbgPhRFXRwuew0oclU
pWMtUyt7sWohD2dPQVgYf8U6enTmhlHzdpEGUjbm2X2hLuSDjqmKDaMZB3/OG2n/uGIwP1j29WVg
TOGX84uOkimvBmz84AO682MMbk6Ap9Fjb5JGuxRUogK6NbZJwEzh4JzV9dZIyO48X+ZQ6wqlP+0w
Z8GOHRnYJwLFs5ZbE8SxN7PI0Z5tP/sckk+fRcLTJVqbz4i+GJO15+mf8mdt+YCjT2dgcMa3SVHL
ixaKsmjkfk5UdU/IXYE5t2/dL0M7LP8CQr5IS7mQy9/LyP+uf4FjvRo/k3TQw2cUsCmdFFFyL0+E
D68/Kvgsc8qage6NQdvfv8KJr5HfNd1YB5WKdiC8ws+/uOYYrH0tez2VwLsOj8BCzVLS6LI4Zh7L
c6rXBuj5Z6HN+2FsR4HPXVL/14l5k/KLa5TfVnWdoqZV5k//RcxpDtMQ85ZeDvY5osojhotOo+nS
Lok/vXgwf5mwIi0pA9+GLtawC2M8VgJgfdO6AwCf718X7tGlcAmSAiqQmQo1db6zEM8cZxXGZeEB
E6aXP1M3xWyTPAFnUKikn6Iu7cXGF4V9VcHhky1RkQBIsL3Z/0CRBS89TrAnhlMO6qoE+1sVGEMo
c0KMtv9MXdfpaow8YQ73p8xpQ+FunBE5d9F1pELQ14OgV+FqWv/9GeGWcxssEBGgo/D8SHUXC4wE
DaoEgf9iqosRzCSNLAw4FNqM9LPTSuumeNWW/XHw0XRreUxyVf5LkfB3r2nfoVOi7vr2y2iUvBOD
HrmXjM1L1EuTMIuoK9cvjlM7mWrZxvQwFZSwAcPY9jSlgXdsuwHzJCoJGibOhE8TLDee2PM+wO1y
ii9TYujWVCJ/vAFrB/fZBG7vrILo4pNRvg7KvEvF2TOuE2b0wVMtPvI8Z/QNzu9vV5useInU6fRA
y/Xg5IzfZHK8coCg520GvJDZiBKRpYUXV/R2Na5SAaKZNbMWWBKD3H5JoqsUYTlbiEhFtIimPSqr
dE63Y6BW/8Tb3iIjFuZ7GgER12Hiq0ilrH7Vl3qgvwpIp6EivWsZZMwGg3spLFO7MI9rR+5sKC/z
8VR4FGdezpSIdczzRbbYZdQfRMYKqKS9Gr4h1pfIl3+23Z/jitWQ5RwJRrTMcbCEoge7+Z4zVQkj
B4x48fka9VaJx6wYCF8ZcrjXFgdfgB5VdodO6UTSBnVD9yRsiLcCNNVnYCIEOn5IOHglVfxTyat6
SnDxZfGgOEhJ/69kt37Im68DRzgPmJRde0a1si3QoRlMew56gsuMbv9HiTn/bDRAiyUek79b9+bh
3D07QpzgCPBJpmZlME3tHeufg2ZetR6nLwQfq/TO6k0DWKGA/ehN8roO/5cUazhFM18SIRXOQ58Y
CyIuDDlaY+tgOcKNf2dMw6pb6LDDpBJJdDKzf0ay7Vy/fPIQ868VgQkWEiBPMOpRWuDwSDWigZLJ
IJVyUE3atfV65tO3KIGaAFDRn5B3f4lkFRUVWo7ERV7q70WVJ2AxM8T9bCX6XrRZSBE1dBfoSNkU
eUBTUIpYbGjo1qkIj2tkD6LJbGoVG67zn68SbMcj7bcF6MTbSk4C3gWoazU/iKaalr8REAAcsuAZ
sKYW1lgxkgtdAGdXshu/WmrFZfluIvYr2QNbOklqFVkgg6kDSlOeDjXI2pBDGC9OyCEipWJ3t9NW
qKeYJzeJoOWsdVHBnlftml6UL4yuglG7SmgHWHg2artaUpMJ9vH1CeruV6hE0Pc3NR/ktXCgqy+x
Lt8ILvAoLGmh88CSi2IVVuOTNqvXWSYDsNr9pVksL2sTD/e+V3q/COxlHu0Wym2+sEdUQ5esXKup
nUrrdM96IxSaILozGFWAniVa4zIeQHmRpfOYH5F8KatfWpTTnk/RSs763qM9mZdFMeO6ESasXIE2
5FM8MeQKhSGaLvpJmEHbDp2qim2gUE3OO4g1pKBvSjJiUjJxqsfJO6x0bbVsq/N/r1ITLrEL/O8Z
1NKrfFa0hqskeY7waq2nJ47pdvcyow2+8j1vTPvr9CbZt2hqfiBTj+e3KD55NvCmcdyWVJGBiAKG
obfz9GO3CsERfTwbX+EYtcX5x8PRrQ+87IpjfprG8JXrARushYT4AGcJlUQxn/+tuQjfEDwpCzgn
xAmkIxB/NXUzKIxaSA1Tf9jTA/2+ZYbN0WX14gALqjvfw3s05eb0o3g2fXmIv2kAJ4z601kHxvq5
xZQOSRfP+gaYdAIzajssaVL5xq8y1UDt2BR1uiDR1NKsEksNWt23fFPniDp3ZPoenQ651/zgFlJo
vtMLC/5q4430Lp9ykS4xyEsZ19vcPKhRfzX0O2oNvQWH0VfzxPN4A44u1mp7BhkHZG3rQBWuPTjD
2hjcHLS+b6VkgvR4o2L5TDf1zfpXH3PlVm6Rw3P/yFD/JFw1MsBHhUQsjutiixVbTammX62yyP8r
j0cEvW3zqKRDzoitZYKFGlQKJwy5cV03nw9FK598d9qCFeknF/AC3/N42d6W8ePH1VfQtlq4f9GT
eJPbj1ZAJbfxD22aQjbq/nZia5mc9CdWcjp9cxs0n+RZr7gnmT0SBtqEr3iErfqFf47NYoDGKe2Z
im5U4cmzEdgGMlJNcbNPpKxQt1G2KBngu/rHyDZjhDKu1ZmvMIvYzUwhnEjvB1ZEMjsurd89lfvn
M6zlmUo7sA+3vzCrZNJtQf4UtSi1bz9QYcdZnrIW4mLMBY6IRZcX3Sl1J/n2AQIZbyBwzAZwh37B
iVmLFxkiIJ3fRjeqQen3lCB3Us5o+jSUrrbWLBGr0AoVnDGDvfpDA6UbCozIByRiSaPm7nSlQsuh
soj3yX7X1qthxOT+K8uDQiSK+ADHzbmuDP9ZPYtQq4L84c0BjKdPQb/l1xQgYnTXKGRrAfCX+Xdn
hQx3x1cKtzMJPmz4Anbo+BSHhRIyxOY5SHzcy6XjtQ6K2AKPliT6BqL/uBxiPJvqH+piRJQkUzCG
qZBMTw9Mru9MH8urwfgGtYH7BwbjjA3wuOW05flu1wUuCbZVzeqS7AxkrNQzi30sIbzF0capk4io
kDSRw+uHfefGo2XY/8sg5TM1U7odN1pFgpLgPFUIkGdwt009vJhpORRCW3LySJJ9ZtaN13z/FidK
mD5D5EcB2k0NEtEbmluIOWdtI5QJxvddct6vAKldVIyaomtBMyG5e5X8UCv40qtHM/o2aQCXbQo3
xH3hAZVIj8O/sheQxpb6llnpD3KF2SEB57SipJ+IsvUhquJOGq3FZIHRcmFKNT+FtLhE9QBJhYt6
7MBOx5fbRNj89/iJ3sZslkXR45XQ9LidCTPHGj5ujETlnusHRsMQx8rpChV8ZeRLwN52xzKMN7eU
Q0uVRMs/5tBiOMZAMXldnzDpHxXgFiPxXQjpCEIZ8KTD4HgS2JuZljgSBIcZ8BjOW/5QwLpU1nBC
SwIuPm2frJfWikKc7ztHQpbZACpWD5GTJ8tB8e4bFdPKThp0nihWHipqmF1x+M+/zA17fhLwoVLP
40TR69dadbHqAUKaXbNqCBYyl2dIkspFoV4pCWBTnA0h8Ctrv73L841CTq1GSWcty/MVur+7NfA7
Qa2k8EiNYHlVK/MNZtRZHF5UtOly/7ix774soyGGwjHiWh6vWQNTTH54C8dA/vUIixLR+DBm5fec
/w+tcOiUOmLTb5BcP+WVte+O9uVVH4aMctZBirRbZwYcOP6QRIHBht4NEC09jtCVtZ1em1VT86ak
16nuCXESBxkYbWF/djbWMVCHqL3e0dBu5pDkscpi1zN/BgRptIIpw9eQc5WFLrAuUijE0GD0w4oi
DelkWbbY+DWDgSScZAkdE+K5KW8Yz4/pjz71+4VhHlYP+5D9xv9rvinLcW/TAaxFr31qnmHbvxVg
Uf5aJxHnjDJ1TyhWJGTcm2dKraIFW/g9CVYf3SHoirSer/aqPV8lvnHV36dZZ8BoSteM+0KhLvlf
uKeyE1HMwZh1B3QDh6OG7hpF/Pn4ENtR9llre7cnYcu3FiWfvgjKDAzHmjqYlFInjRb3KImZLM0q
4eckuoy1TnjWLSEG7Ui1EnxJqxqmKxymZJ9Ze7CUs5cAB2u9gClw+SGhhXfjtLPMPGnmsPbkzFJO
a0zhkzCd7ylCb0Nji6YoaElHsfea+32usuMJCSTxdiKZZe7GkO0LmK/AmTUtWfw7sTS9Q1WzKj9y
4SC0Lfl8GRpPPt7PkS8ftwgohC6++1cszdBA1qW6ivjTeyRNKmbiFZ8pO2gLYb2s4r1vovgBS0bQ
tnmIK3AIog/2uQjwNmN0hF8J3IfSyeQMJ72CCKtPMKJWfiFPWQkkWlYfosbL8JVmv0RTTzahJUSN
iBNKLxDq65alQRW5llMeEv9Td4TyVdicdUsVJfLq1qiWlzLHAuAnKpYAbsLm9j2XKTFw4MweZolB
D7pDuAoY3Tt17pTMITVMHQsmy1KmQ2zspGbdagpkwptHHRJsxMOBjbiCzAw9nFuneqrDbCOQU8NX
rfXZjokWX1dVryf1cBJm0fc+n2Gl7JVsGX2CdCogQM+UTphVrGB3/O4ZNpZkUgU68UpGOCfn/Kke
W5tOgS45zSln8qa0JJ+jYhIPSdiSOVTqNLcx/kv9J4aQrJsOIsDkdxFnNbTWS3g+9z3qNKWMVvgx
VbfV6c0N3TWFbSI+tu1sXMIFYLGP2COqgGFVckWB4x8tdMnYUdQYRTtuz9D3r7V7RQF0kmzerbD+
DHWOh+0GdfVue2g/jIkN22w512xRw37+XhuiNsGny/qJgZu94ahPjxaTvoqXoJ5s9aCphYLM1MHV
fOV8myF/M+C/HgKZ4Nw4GbNP6dAmjhTTh5QyVJosc1uvsbdDEhQOdRvBFchCwThoEpZ/D7lBNS/b
nkex83oRCQr52aEPE+zTf5RrECJKf3mKgqF+4SrB/SnrFaBdLuXI954/vGO5AMBiO/uj+n19zHBc
OOC4V29ouyAa4TIp1FRdWSrNkKVrvSdKK5YzhGgKqfPDUhP657p3mW6mraKc2WBwkvZnwGUkhu5n
m556A1hIDCc8ITSWdPBw2briaA5BAZ6XxE9Dyd6nJNCb3UiZiK4tpauntDRzIJoxcXQeZ70O5r7l
AMfL+z4YF10n12mvZD0rOQ9Ejcqwpp6sCGSvd0oA0UpoZYOm9e1ojnG3nDygBj4X1GwZpte3dI+D
5EqP/51HkfxCwP7D8kNf5VBfYJEe3Fq0TeGhPAiA6az6nkPraM9/Er4px0oApclGQEJWUG2sujY5
/vA/t1WFv7gEmkDb29XEeiZuW7olbp2LBfhIDNmbOkfigFpBy/Eo8fH6mXL8bZPzIWjIIjGDJvtI
GH8wf3ZS6h7MSTwGz2NnsNg9siMgP2ILyuA1J3dbpGxOhpyjePiMDVpiLyM/p5Qzi5qubCS1kShQ
rmT+MVu+i+sp95p8Q6Qw5qQS6yleX2FqTj3CTJskyFwTexdtjS41bVKrtSjej1/s1vQdvOzVbg/O
02CgWbwXD3Nc3ecRrliiU2b1ZcMe+6ESYNpd35bqG6YHW3BsvHECGNYteMY63p7Z7IeEjf3PahDm
WCWaSgj20HOWivyizV8LFM10uY8sVEcaUd7Inpf9eFcH08KJYLF2GNMjWu/mExK+CoT/SSQeHHl9
aatqNAO7cgy5W1hwPpR6M176s6wazp36f3CMqDXxVPctCA5GqDFoKVB7GAyhzsHllwHmMuodiCKQ
65hJX5jNMO56hH1OgNZEslTssgzZLtVf6vIT/x7yx5aiYaYw8+r7+fTk6v/9uR9cUhBhjDc8Ic51
FTzboiuk4s2zZ9xscp6t2zadesIND7/ncRemKjBDOYetsDlCjLwgTyVnkq6ofV9HPh4zwckv9/KM
01TjVf804sqUFaz5df/RWAusN3R5pty2h16BOfd/khxXsqbnGuLoBp7lNP/tyQPGKE0FyQbbU83Q
BC4QK2lEaTIhCFYvgJZ83ypGcTAs2g4FrD5++uin8E81q4HGczr5AqJ9hH3+eMP4TKSqGTPqSZzB
v1SPStd4U1AJS39/UJUIjb30iNQkmVS4xUy6te5RdM/71RoLj+kEe5XokYVgrx85Yw8H0F/cYJyO
UhfumARDdSsRnanMKww+FfbTPDknjPRpophuEOZiWLecpC+vT9if2moyD+LlC4o5w2pOjdcqGsgj
zRMRWJ2c0KvGFkRgvMpHagA9fLdmVSjShgYsxFATrsQREoiqtO103H19LFPDFWnUexmDDChCGich
NyGnhLwlrGS45B76zQyzw7bflFdZDe7x3M7UWkqg0V18aWEGLJnrzXYGv35RuMRhB/kdk3tt5hd7
K/vUeIvSfkPt8ZNdvJQo9o2nUJQ0b/7Qf5shQRSbe6sfYn9MGOAjhr8IQB6ANmwJHLEwKJYcVasF
l6tg/MxEyPwCV24xjx30ev9ynHdrPRuYwjX4a8/DpoMWYhQFMqO4mBCGfyaIQcRCYLAY0K7TU5W/
WKiYoEaVfJDzqivtb4ikJ5Hw/iOV7g09PG39b2hYO2acEG97LGXZIv8CnGoejEEb5hHNizn3Hbbq
FqWAEw59UMV9qXyFshcsDW1focCRYkpZz5nsiDXUGxM+6kchlz3vCUDYkz2x5+e3owTmnlZ4JZSN
/juQxxnFLKB/DTyxgnnS14ryGD5BEUv67n4XwHSaCFV0o0HcF6/tJKHr5f+zKU2fl5MGHuUfZ3l5
bh8QpzkYrkHZO1df3Z8XDhG8gYH2Mjo1PMwPWRf0/BkF/NPOFyQtbCsajGSoTznloMUIcKWKON4R
PxvJ5bbGbKrCBmsqsz49dpBjq4Urt/lsF+N3Q6ca+EBwimZ4dsZVm6auCMNB9R3ysjzx7xBJ1XfX
xIIjKKwowDIdU6mx2hEBFFTW5YhYEGxRL0t2ITutvY5eUyk9CXtHtrAmrSyMHiCr5BodCJHhQoZq
labWdr3kvoViOlO6Nzrey3PjNHyGD/q4wdo2N0fYYHBTS8qayzVf8hczLEnpAz8Mk4tGcXXzzmxU
89qz5xTILfQH19L4uayxT84eF3MK8wQsKl0lOyncyONbGuxCujzccpbEhBzUnl3nDXNWdpLMPNYq
0xBDW9dpl+fcmwBC4wyoKyOi7Xm9a+6wZkhZ4Vu5KL9Y2zNOk5qO6MNkhZLrpjH2K2qyc4fC/qIS
FDXnOcrQ6rgeqBfLqiEdQ2pYZb5a47tThx9OoMP5cMjLwUpFFh41sACzoJ4kvwrdcNBWHRq3Owuv
xXVFYtCseTKiAB1VDcI6ucZx+A5LVtFOcF5r0Jf3k9WrStLlJjy+Wogu5w7xk5h9WSrn4IVoQR97
5VUov1aHQ7AlT/M5lAk1ChSykv87IrF7WN3EiWBXY65bYpvfd4JP3ddSby9u6dWm6crhJp13flZ4
PlPN3oHaB1x7bVAYlNedqtQKMx8zVF6SUZMkQKUcDV36fwVxb6Nu6eT07b3maE5JZyHLqZj2Fzo6
w59zdWfdXfAi2v3CPKtlg6cO4leCAm2ceCyC6tIs/jC8Gdnh/oI0z9KE3CtQMn4nCC5Z8u4vOXGi
ISrHe0Re2LgFANbwMrcCroZUru5ioyZQtmsDckBwJqg3G1n2/mkYdkWZwTW9VmQc5I1gxZHVZN5S
g57Wi+fwKqeR4pYP41c/MNV1Hz32qhCD1nh0ADr1ysgt4Dpf9T2IinxmkbC5Eik8X5tttWtknhVq
GbQNmIj91Wt7jTA57VQSEdSmTt65iEbhkVYUVMA5dbacN0vwOXMAPy3whaD4/SZ4BAglE82xxOOM
0U9+bUzcpeQXhni2M9mYlFJf5utOsaab2U7BmjMPcuSxGgL3Uaxb42hQspyalPP9NTxddZ2x5sCz
Bx4aKT6T0LQ6huq35Drblq9CY4FupdvWcLcchWbsKaEBHBDrm8xeOh8zY3VYzOiBKI4nm52mgi+V
7Zau2tK/bKo7Q0iW4/Nd8/McO6KzS1+fCaZBpRd9b5n+J78GN40ZVOq5SqK2ynlgrOuyDIK8OZ5/
gtusQ/2DeewNdWx0utjYToCxWT9M7sGpHTpDEUk94RKY3YGSQ4HG6i9y9OgO8SKJO2iplZdU3zuI
VV/8+FEvwqTkzG8mg7HZdEbcPOuDa1A/aaUN1KhhGSXgtPCzNGFMgf0hAPxv4mJf3jDfFV3ESkg5
b2HncPX11UsQhT1KDhanOaOOYJib7vt9wmgi5coBPrG67pToQlRJUVoJYL/546XDcrf427hfALXu
EZ6lVIzMAOUB7o+bB+Bcy6wSa0/YC53WkNoABox9/zEIMigvgJz1Q0DTmKw94p9azWcRRpZqQnM/
vG0aGnUUZ1ri8YpUcjdMSPmy6tPnNeRwfZuMbZnjmpdGP5tNYaIYifvuJzBY5R8gqEqud0+DRQxp
0alTmjYXXWaKjD0FTaOJbl+ZRFnlcmLBToTHi5tlVXzOkqEHdz05NJNPcP7EFPB9PpcmTgeGh5kf
eADkryo8c7Pn3frG0I5dDuim/f1AZpRyrkRa+yOPJzEu3JEno3uNFEjQZhuIYmqepZx6Oa3sy+Dr
gQgxM9IlJGqPWgpzIqHB2E+whrI8k2qthq9o8d1ic2Ekd2muY0TenGK6bA/qUcfR4s9H3Vjt+rPs
P/DyuAdF95J04bmGlvTohx9U1SsF7QjqsBlf5DcgZHPpJGxsd7Qik98E+Fgr5qMckc07rdNqvRQP
af8sAq4zSvxQWrVkgTa6+BKfqDtV5tfojKxJk8rIH6a3+hEDyG2uRswpz/HSM8mVnHGHXlyqPv7b
nOSh6ozEBN17AWY3Nt11IULSFMrdU9saTmb8RJNaz+hnaONN7NROHTl+V0IbhyutNoKSSrxREqzd
4TvvfFpTaqHm+d9eO4eV5cwbvwnysQdny2SpuvgxSXQgc8Swe2eHLBDLCFWf66hBlUzmxNhACMvu
451J1gAlkf6NnVX+Ywjnxa1CERYqVuU+HuXl+J7ng9Jy4UVWj8OZdiQ9QEiBelUqTev1NTWY3Ctp
dah+ib9Iuj6iA/LlWeELKg722TzlpAxpzfV9zYM8JaRafsoiXzWTQVEl/lm+5v2MPQwsKp3s9RQP
HAHeCBvfANhK4C8IEUM99kL7CDby16G5X8032BfBkYbgd8wMZFEiuxnZbekSTewohbxk1dPhJMJN
3tlVeOVLbk0ExBo93of65MujofNFg21VY9nrSjRfR8Aj6lyH1DbGXXVEbT8LlKTxaXwMFxMVU1Uk
9pgVOGeiXJQG4OT39FbDb0Xcftoxm/erq50kpPD1AkSOcS7MF/76l+atJRAyfrkV8CPIsUHvyFf5
9D+X+xRK57HMtdbGN/xsA6K8TEZqOkFbCj462Kj6C+UXCc8ARvg1zhGVXYODX+3/iLNDsVIhQMu4
NFFa4xHXmaXOuErg2I8jwNY3nGob/4IcNNufEEwxEJkbhc5746667NIAlmAW8rQharPz6gtG52UW
RRQWEp+MUYfJTPhEa410IN4njr2+mj3thdNS1uBdq+q+yoogrRQXaG3TqpWOH5GYbYeF+siVlRqQ
mgDtfcDW4tTWPyR/WYK9RfGBhx3tVN8O7yfDWJ0wMWo9nM7B+f1pacY2VjOnv2bQGfmT1RTm9hjW
t7bPsRAbaOWk5nZDCOUS0uuwSY/D/OAs9kjpuSAeGGBcdhMUhfR2wBhQyOodFSvKwmJCVFPelzWb
27gAedQfheEcFc17uqoilHjTsYuFpqmJzZZyA16YkIG2iaJ4YQA6YulRr01t9y0+FlSUzxOpq+z7
x2iKN3pSmy3VgrO1cyC/K5oB+mBHBEzqrItV90GnPiABK6OcjdyeoLhqLCGrnbTTdkKqJ/d5wQU+
FWc2mnPdG3C/sH1i4bO1NGZ8roplJIARVwRBWYyleMyoRWe7IuxXWNT7X+0cSi1AtcCWhVWq7Sjn
wSbtQyxr4ks3u72q4VvvQvnKInrLXmLbJnqThSQKlOHvJE7CPd8xvP0bVXTxuCELCgsQU4gdQW6S
3EklcxUMpLUt5AtT9OiI/VjbcIcIOnRbVQmwXVDJpUzPYHPmOsNHp83cgy9dpv3i9FVHeVM/IHoF
cTuKUMyOJM3R6BUPmv04UHP/XCOLolHX2vmD20D7RGqgVJsvq87VzpJzR13oToIPIoli156F0VJM
UlRGySZzg7o4T/8g0sVnYV6HJD4xRK5llTKDd+/rHM+dJrfm5DjvxblGvMmjf8CYGdHfnduLC3pp
1hGNmK2zO17RIO41DWaDM7MFyPhJltUX++dev7KaX6DgDvkVJkDH0cXNY0z/xeR78ZKMl9eBdtzk
4aYriqTtKM1DzQ04uNexjtdyZQNtOjOjpc6GogDKzsHKngVh7/gxAvIVzzDw3iDo+XWqJfkhYAe0
p/C+JlNNZ3/wG6V0izQLJZi5UpeYm4MhBM0fSw95K9LZt1MgpXF6l9falWZKKOl0FHwzTHinl3we
A54kicZwjBHvqG1JOApA2hdSOFRplioEQHhN2n5APTu7aB4USJXwrO2CleKW2zLaWIDhqCQXeRSI
Icv4/MWRbFYMDVQm4JvvLG5ix1cbc03+MRZkoD7WcWc68+ZydO0wJIZzNACB9J+MLFeXcsKLdqGl
zviPMQEAjeVk87dadN8NFNBpN/1N3V6wLvRUlMr5HdXaZ3RM/pb079s/XrXweQKxx86itG/DdAo0
/RaFuXuAHLYEPhqXZlNfAC6zta6UgwnXnbojC100N9ej4AAxawlXeiMfqRo8OOpbuhRRdwXAKcsv
C7vgW6Z7AjybpshjS5Iml1XMMbc9ROA8CT1EAY40ztEiMOhiP1JK6Q3ZtQwtyHcuDqFq5oo1XIxX
HZ0rxihmbkNYa1O5XyP8yOH8c3jRllTgARdyH+dpm1LqbMMHe/jPQLne6mEuJbBhBqWqse4H2NzG
CWrGejuUtFJrIq94FDAS6KpGr0PQUqXk9tek/6Rp65We+pvccEfgcmu0kd8nf4Ncsz9AKOxOC1ns
uaF5B1qjr0N9Adnr8AnQbKtaKqtEicw/QeZ4t7RVxp/SbdTam2OqXtbNDz+wz9lZpI2owmguiNJT
2uh5GM8btMBL95+ZrhL7KkYH0ElGFbbF2DSPX44Ftc0Aw2PORJnDaLHMbRHZG7Wm9oqb+ylC+8E0
A4CB2o3kg4JX7COH+4Uq+HtpHPxF7BHTWcQyh+4w7RgBKkjpqE5AfTBxZkpLX5FYBGGJkYLkR1g3
YZxav/SN6O4SGmxKXLFjEUDIGMbDAVG+bWSAABWah4ovN6lZd0/+TILBGwlP7+UrBIziE4x7VB/l
BCV2lHwdf0I3lS6NW3sJWhG19AqJoseFTJ6kcUPYc6R4JWa7WNR1YbFknnf2xlylnYE77xIIa453
5ic9AxbfC0UhWu2JT9pRmXvhty/6PRz100aVtBS9TjbVC7O3Kaa85Ek7xwVTOoRs7x8u+/8SY3k/
6+7LYWXdkObKyTwFWsfui9Ymbo8RM2Txcp5nHUwOqh67mBDkfXLOwLNsZE+SmW9jX8ks/zrjwCTG
z9mSL4AHQDZuZ6Hnj3B60NvCWWpyjD+FlOfRjMwYPui12vEcBKUE0xfnrkxAzeg8cLk1VLhqlhFq
NUbWggnQhHFNTnQ5uzY6+tS5NIcBlISJi7y/9owcyc8deTTIWDGVjvfwSHGh4Pzldwd+ZZa425/0
9+W3GwJqr/znri2YjGoB8pYxVpYzInvZWKzk/XbmKZq2eze5LanmfjCbYoPXybSU+EbofRKJdg5w
/kbViws2muEnk3M6kckSvMankvlhsWJDdlc3+e+azT1K9XukxhWlksK/CaENTCyZf2XffSuK8I13
pA5aqxMD/JBwKKNdRoRa0es7+Xjk2RdrQ9HvQvNQ2g2olbZqP3JkZgFRg3pMf4D1tmuOdXdTcaAf
LHzadsn0YiXzXj7LNxpLiqvEp2v7W5HloTkRtsJm+hg1uh8sHpsZQ7bOKuChyyuq0adqhz+dh4mH
GIWdgMg0PICWV5H4wytlzU7vN496yRY7ev/1OF2KQYXEJQ/s7m1tbLgKPKdvoIoTvxwamBvP3SyV
Etc0+K2r14bmywFKDD48r3qhc12sXh8nf2P7VMXxN4dFvx8+7GGaYe5GRw9o1Ue4Y4Y9YbZ9Peod
UCbKfaRP31+aiyONOyNERWjyPw9UJgqaW17ECYcypSnTXxct6NsvrTOq+FHHt0SXJsi6g9FiA4B7
tPOO/zX+anguw5pS4Rw6XKlxOy/HwfTppbfC5y+LdjE+MApjfWLJmNIdZ/Jylwt9HfvbhxjxhotW
TwPfq+tIZhOkSBgDgzzYpTD5lZfPe6r06AL+bIqCrEuc22FUgtm9PwkIrWNvMWUZCSEMPdrosTXv
XKGxxcKIKUr5sSPVypgmDvqKGd+D+1Ib3fj4jE0OoJ4OcJmvq6tgtf35amlCftURg4NNW7o/Bw6y
aO5FgmQSRYDIbeTZ+/owlZRjPiakLoOCvrgCGALxQRkPr3bqra/nxzr2wtuxzG90uVfZoJ4S4IM0
+/NHtant9bWbp41NQNVqsuvy5nHF0THPehTKn5uAYeN+icvbs9jLL+Vyb+J0B7GLb7Mzc2I0sL1a
NMjznbrtYsBnDaZk4qLJhVu4LqzJ4GtSFCky020L1FucuP46Dm/u2ntMjOevkRJYXNxPDG5IyCgY
CfIfR/vltE9KfBUhYYv+DS+tWQC9c3cxEDRqtww/W8s1c4VPNlDVPGo4P78qT31xq0nNxWqrOH72
ZCEyzEemAeptQqyxP6lrjgs60Js23EonuM6B6d+bNHHVBvdrcsBmbTSFZ8f6sAdfEOrOHtm/gHOA
E1U/Vq1bT6Uuzb1cuIi2yoL0rnQdLhqS2g9YXHBB4+FlDt8mAKtgrH2yFKI5/aFNoAXJ81uZjaFd
TzVbsjJA2fxsm0UbNYtT0pooycM+Aby1lPIyhtfatgaVa3aT6YKYA9By80o2EIdWeXmk/AWVZCqa
OxcHegdoQk97XgB5gHNy/gvD0FAxBm9fyV9jy6joFfXzByou2J1L66dvj+04iMu2jrqX4E+lP368
CTtGf52EMotIMjxDNIx7C8YmQtGlhn1R7UtLMlQB4snLfgBHi4xyIZ3u6R43Yks1nUbZrPCStBHZ
Dki4LwxIsR5uvTmx+Dgi9sli5opB6MnzRTta9DF5eKdPrnrYmKlHnVfcJrKJBS+uWBs0VKGnIjw7
7p8JUQxP9JkiwyYyq4KVWeaVIadNlFyweempZFrEdxVvpacYoBb2RCkwRaBjYK4AGTIdrYDC6h1a
1Hb5O5ncVPUVIOaWf9EuAo5XDLzIp+fBjKY6mZTd05uMa5qlZ6ICdDxFveYhdcKqpd1zzEhOhf0C
5zPS64FHbtjn8pRXSR6/s13dO2S0/Rh30hP00gNtspOiUr9rJIQcRLIivq4qaici5bZRpIJFyBhz
Zpxp13MwrCbmSYAfPTUiyb++23Oq0b6fSn1F8HlhPGSQaZHkCEegF6liI93A6ar3nYcnOWAOwDsx
r2dDeiHC4f2XvmFZM1LUzCY4G2LVLZ0Jbq4VhhTBH6YD/AfU4bF2oIRGWijssInKJ56lJZAAYfvi
Yg2KfN2GeTTNWCi98X1eoUKY+rezESTRp9qgU8QFX5H+zPTuKdl+45zY5XoPlCYicEXjrcKpwS50
6QdbzUhKDcl4L9/eLh6SfHbbI2U7xxtpCZ0Uly0EFZMRSI0w/AhL1yG4YcLZYUGCuT7683zk4Zpw
gC2pmHX0NxkkhidHZ4bfM71gPJJDs4xzaL1E0nDHaZSP8fJEYOY8z5CkpZUwUB5uyNkkY3Yibfe8
x7qGiTmLIxO7SrpizEZDWyiOrh4SJ8e2hOl1gW0eWGCm5XLkVEmH/UtBCgAYChReMO4/TEceEQFl
DxX76FAzf7K5q35Nl5who+04JFTf6wu5rHJu0Y8koayEsUjWHzYiM2dL4v0bkVQfHuEpzYyHFWdg
ROYmERmRaOBHavVpHw6juZM7IQowCn22lHFOUSoDxL/ggljCcUvA/1AgtnTEXxpVRnd8md+T14RE
gW9TvjHpsyeZ3NWu93U5Xoh5AojgDIhtZKkX/eIWZbnXVM3uusoGHiUHHS2AUAl5YvrH387KLkIW
dc5J0/9w/ZBWu1fcjMThTQCCC9vQNKuzmFN23ZVjHZ4pgJmY4og+XwmEpAmQpUD/OtXvHW5pj3WC
vJ1J9BDS0WzFi7LD/drWsfV8SN6fgVoE47w8Tn2rISdsRZaF05W3cRbqjUw55YwIMyHoT9s4lfKN
chE0l3cHnJkLjz/40AmaxVbADg7oCh6ceOqZOZMQSQy49pPaZQLfBCQ5Ujkz4eSxckcZr3q9hmxw
SPPtNPWKZgiLeFr9QYvnuYT86TXnhhytSxpNw9jIh2ABrkDnLvfDZACv5fKlOMx4KMmAyw0ak+gE
JFEy1ryFaxxUr59Rk8DfDdP318GoC0YpCNxf6/UpQq+h2tD/0BkBXLJDHbvF6T8vTLOfuvBKkybu
NDzL3P/SxDjxtEH6tmS7vmEyZZRvW3O3XMWU/narwIjf3a/trhmcxwf1dMMmCP7tY4xSF9ZjxTiH
L1bwt9dABIjQ6NcskBZ6mw4GEl1Hi3ubGKXkX4fb0B2hv7tGg+Oa2V5ttXxCHgmdgGLz6VotiCSt
tODt1e9n1CSFaVPCFZH0msXduudf/X4aIzkZ73IOkSqo8vuITHKIs5vGJ/fqd4qrzjJrs4r7oz3r
THK2f17xfAprCqDpUhZxrAOVaQh57mEZweMpdFJWMIEbziCkchhbJBbWYTL62uPgUDV5l1RlLTVp
myCkPTQ7o5UyJCH9QvTbrILHS527u2pO8GcxDKmOe/TkHPJjFO93YFyRKTUtMStiixNXc/tK+dnU
c2MRQHTgtHEliI4ppIaBj7xMwswDD7NQSyppObvGC5END9t2lAtoyC2LVL7VVymZuZ2XCcEtN24+
KHRJSKkVmRkOr3A6Yg81v5JLPsxkkOQK5g7mqrmg44cU3NZwC1aYY52IL2ZajDBPjXAPpKOo1ogt
g30aUD7bqLNhoT/LiB7fLVX6XAh57wavn7x0V7rFrCH9HKlYTiU0hsEH1D4YBIplxC1bBAvIIdsW
p2zDi9hvKKenIG51TL25zp+EV7WxZJxg2i2qd8D4a48wnrKf3O2f3MQMjitTG5HiOTdkQPj1d7oA
iXA0zlVEBmoPBTEgMQBPGkxksZcvhPmVZcUUrpFKePSFcBVoHcfyd+ydY3guAM6doGKAvMNURgam
njkepL2bf9Jv4v6xKU/QWITm5fnfxs/2nCJP1KuaaPQ9NapVuQAsLdijo2gZFfXCkjvPdC50p4Au
LvOQ04Uj84AIUCnVeY6GpeWhuYbDBAwLFLB7xUneeKz3wSbAm8HSzb1ddtk1ci8+blrT/DiT7wdF
Ci6qwkRrF/7nU5MJl2r1a1+xlnnFGGpPv91ZmqM09SHe2Z7RPdCRHFVXtRCCOn2k9TlE6+Dw7nop
EMLm3SqdKG2rHxqlVFbV5zAMBoIarS+VN+Rk7wYgRMGbLZCA8tGgiVeVQKOQbb+HSnIdU33BhFef
haBD2bBOlpNxAWYPrApqjPurNqknYKGhZe1MpnXdW6mb8xQQHyBSSus2MeTkQbkdRbhs9kWIaFtD
nN6IFhq2dzWzwjgNp6ICKF0LluPEQ0KUIzxws5tQqO4lJkXJKlrafyGkYQmUthuEvTOC6GzP4jWo
eRFjZbLKcNrUIZRhBhfko+qlZEzqqAC/sEGzKe3M4Vrlw3dQsRZItEOnSUoQajtTT4AMi8axJkVZ
mvqYsTwtStjOgyCyNA8EH0R7I5SSJ7FbKgoHuR1lziqXTI7Yberxy5rpGcaeHVJY4ed2kiWkAB8h
aqh82XFjBpfC6Qm6VRmByz1ekxIIV1AQ2fA+d9vzuDjeyTYYCyFYmbT8mZKuHoa+QYUa/IB3M1Cg
9uq36c/IrRYFWCg5wFeckx1RmMg52mIdnOm27v/LWk2lJcQrP8ud6imbLDJt1VA/b0VT9OFUODPJ
0qrVPjSqI0hMzMTtQTaUZOFipDw+0yTHumT+zJN837/JhOXG87+EymRZqkE3+5uuHN7hsVjJQF4W
OH7blN4RWccd4d8ZxQXJaTM9DhcvucsTFmNGPVn7iRynxd7FlEtAp/Jg0pfUZ6ufL3iwmN1WIOqF
LrNCRiVCnHlmijvwB97/ybwTSbGcp6/5b7YxFHyRMMnbWXY41LSS/vj9/GGScLSgeXLEvvt3QgAq
jLXxDs6Lop3gl314QaqjzvA9Exla8oZmGR4vlBfPJBthMjyHVYw6rYuzIrSVHaN6IM0da6OTqSwV
wNRtZzZDfKqWMW/BFG5Vntq9lmbj4eLFGb5tMu/B/W/Htq6S36ficG6rfLqqsL3nePxMFV/hxBRy
6XyijeRr80t6LecLgv2exjGpyy4oraJJEsDcgIaUxVUFFgcgMDx35VPwoo99B0NBCIqduR4IUqOx
hdjH5iQBIXYhK6897al3mVKTicXl3Y79nOG4RoI6lJ3eGnb/nSXfM6a1eMMZIIvNmlpiNBuClJjK
5PKCop907ltkdBbe4VlK+FfQRYMvfkKK2ngUeoxYHXBTDd/A19/zjKARg2vGTxjcxZDVgHNdsab5
GRdLFARPPv3PBDfMnkCvc2xVtTwI2gL2b3TsLK0+7jK6smBKv/yTqfeAVoVHBYLT1g7YEHUwREkP
mmFeQubnxmel+8yb0vosbj+4mshG5zmHArQ3k8RIzZTRSvWc/NJNFEfzUVWH9klzUxKOPsjS2uXb
51NPMspTMS/Mw3MT3x3txKmNQt0x4PVOFe1fvfX6BmGe7G9GXwVKYR/rtRHKuJQn1FZe2srfK1st
HiqF4n08dX89zdxShkLVwvqHC9newfR6+49ZRUXjrUt8eqc430h8DEmnCMPsAE6YxtFr2Xsln5SQ
VHh8I9Aor95rTIuw7VsqPrAhPNjefQCgMolXQCgXb6rh6fdTiAAddhQQqYn41fmk+EUZWLVN+rOj
rHxocedPg5PSG02u+0q5f/OKsXMxIMenddQwUtcrmjstRNt/yZ718OGhZrcwjl4apxNXV9JxEsjk
HNFmgvoAV76UDg6ZW9leW1f1kV/L+15pCy6QIDHHULgFtWkNRLNqw4ZGyW1B75cZHzHMU+FrkZMH
tcRFcFY3a9zqHzFi9HyW8j/zQDCneTmLa9Q15qq/D2wM6nhUqiQ5cWa6WlX+AVJpaif9PUkuEhDo
cRnApguCFfoSFmIqnRXcYr0UfX8BWTRcB+dqSUyQREj3ubeQf987Xv54yEv2fpPHCIKbCOTzoneN
+jUIhJXnth46NGls5wNnFj1xY/+CstCjMTxY6l5xG3l2FOL8zZq9ZnkdDakFWS4yHof/bfGmGAjP
bTHy/KvhG5COiKKog63IP1yFO6YwpXCzd06CSA4wc21MzqGBXS6JzCtmm37QYUbiDM/MNiE8C+YM
pn3LM3F3NT7ZQJDujSib5Oo+vh84wxKs5qliGKsWuh7K7BAaDyDFxiscuQkgwcS/MTZsHhkodma0
UxeuS4KKjxFLvsU9dgXzx8urftyv8/25hWJC+MGK3Z+/0MQWykhkYnU+Wh7L+WblNNII13mn0CEC
TGeiI+b/rBEdjFYRdtJ8LmoyP5hsfMRHC3DU4HQa3/AsniWOMM66sTyfZH+kTjpU+chRNFbOkCc4
JAjqc8dr5F1ltDmrgCbi/TMOlQA94/kIVR7AhfmhGzAEMc0ALuJPo7PAp2cZr9gfyY16LtkXDfxN
GHwjkVEcZR7b73S13hVX9pdIVSRrFIli0b2N9YFP0lr7neTy6azes7xLOxPCl9QqAwXla/k52zqf
c4EwQ9UBz8ULac+HCfSUpYj6Zgwj65JADeRqJeqHZNzMIUn6tdxwAUm4hfovaA1hRvk9yGLFZVBw
7WPLTKvnIYPQKoxyVuNoCqK7pWfJZ3G3X99CPM7NN/gFh2lvSs52zbtWJG/64AoHTUebeYD4hUMO
keXczXrDbnE4TnwIJW0Tj0dHaHHWW2PNblqg2J42AQeUPAGfYIbqg0kUsmq1UEyE2QJV9IW+oG9n
5QeWq6kVbAbauiesozyZl4SXXOnnp66uXlDLVDP7tbPIUoN7RJVEIWOZNatwlmb2x2JpU/oMR0o9
G83vkzZ4iQkb5UjhyklANaOFg3MX89ajPbxSx96GAkQ+9asFOR46AsMSjYeVehjBgEq+NMWgu3Iv
uNkBGam8i1ctH/P04djbcfTIDXADoEB/8bzOGqQwiAmp2DZeAbGIzR5Qj8TFKveAKt8LqcxbDumI
XzqaYvRNAfSgynrS22rSnii6AftQUhb1c+dsXT/y4jRUiUOB+l/meKP76tujr5onY6Sl+WdftHy+
OAd8k7ZEl7BBJx3oNMassON6Uu4as42ENzrut/O/zBTC2BiUUKYWMDk/jh4B3fgHNr8yvQ7xe9LY
5IpbSjIudr6e+Ecfbbq3l5mXAJXzEQXrVNmkPearRao2NBKKRAM3UR9HZnTd6/yhXyqwLXn4G9Ga
iEpIfj2G0zAVH0/FYM1O4BC9eShjHcfFI0kJ/q801piwxWgzAOCLgEra/o5GkDkdVOJtNtCZ1s7q
WkoOaqY4qNGHf94BW3RiSvmMW7/ucfI3Ph8C4TcVpX9e+mwmNXL7+AKi1pXOo9vExU8oYqBWLTMS
63Ai40jLYjh2tgX1TwTG936YqkbNRaRHixBdd0O8E3NwQHVVziIkWHU4Ke5kLez8gpiWLF8F86im
kpibixFkQvx7dBQGKOVMm6ZIQR6CEAEsWmlkHxwFy68W6WUdlfLlfU0DQBsb2DWJhJBpwMcvf/pG
ah2Ix48IyLUBVqUHXCmuJGt90N8V+fkFPVugljti2SqOwrPUnjG9GiWAxfBSHZf7fmnd4UjuvA9E
Wsm30NXKqc3c/5I7nWg5k+1acExXUmls9GLqM/+ixkqOJgRh4oPrLwP+ktvnza191y2dBq8cvVZr
JkKaHrPV0WPtZeE8NMgqTQN9U2S2/URztqFCW8WtPz93pmVzlxcINcZlK8QUXrH+kjrX77qbQifK
/K2aKYDxpAenjfio5WxMasdK8ijoXDaKBYaiXmJV6kYEBeMXc+QfCX2eSN/bK1SZ94RIOXHXPHdd
csxabQFTHgDzYXorF/YW8XpzWyo/blggFhwCSdx740F38qhQelkF9ZXzG0EJltjGBIneORzbGKmh
fRsXVzRQCWlGaVpSCdl/Or8+nHoKCpJr2A6WbjRzmHpRF46BqksbctUom06k0j2MZzVKxrt1yhO2
3tCPcq3/1Dxz/+ju2vKnnG5bfwmSdR6guMFlwLWAuALCtMSpkvzMVu9MMcG92bXWgEyXpUaFQm7Y
/pwlF33V///v0NUGKvZqElMO0imNSFv8HxWStsHlhsQ4d2fhzuZGqOwsp68/mzSpoX8kgXPkrkax
YLkMRiovaGbWW/AtBVanMRA1/hvm1MlBlaWsjtF6+3hZ4UYLa2cA7QDi2A0yrtN6TLiu7XuXmF0A
lCnKpzOMdDJ50RDKX89K1cT1PtOiWa5A1IM5GeA9zD30DIfgaJ7TN/tw1gsHhR30ia9BxZ/q/wK3
itp2d9LLm/muZ5FmdsvFyqbekHqVX8KN0ZQPNDc6ez+03o0IGGT/Z1FHyfGzrvEEbV7NS9JXpUe4
cZ1+qdWrSMDDbKfUOZs15ErCEZUd3MfahDDxxV4yuyHVr0DKPTSKFgSAWHDy7dvzRHb1CohA66if
2jIhaH6zh/h+fLotKdZqv9s4F5BECH3fIOF7eoTUJuxU/DQIovcjDtg74009QwgOu6SrvzwSeQfK
Kid6xcKfwfBDSZRWRqpq8uVzXUHkuluB9MPCDttLgM6PlVk6FQQAYKHuZgN1JT6/fpWciEqHV8qR
jo/WmlkNBIElYVxZSTf7fO8rZ5KTAASGTEA2tnlOlnJanSxkX0fYD6l75N7bPIsoxJbHxhHEbouC
VyxuB9gwuoA3No61Zk7rDpYRXac7IKPWKRTl+lRTI6JZnL+YvKhsk5M0VrnDYFp6kSvCoK8dId+X
mI+kR2IZAc9C20Hu2fL7kxLsAdRxz4H7sFxhTRk7LCkkaGVV6TfpwXQhhvhdyE3S1h/iecUZMn0P
/oYYrahnFDTmnV4pdzrAazdPuDtUqeteojYCNDCcbAFyvfJD+ZlluHPSt6ddAA6BtGEjBHmyuoLq
Oi91pQJStM9LOWSPmhemxM3oRgCBPhECDF7N/13FMygYdK6HqG/FYG+NGqoptau0DzXy7ilFhe+Y
tTf05Xbem49XVxw/C9R8/0+iEH5wCBvC+8ChZwP1yPQKRZYKWTXW71gouXkPVerlYYEcEmV5D6rA
5RrIESrKny6eHchTWbN7/w5nNbj3cjv8mExWaYfmugt7t3FLLxbtwYdh/AIjyFmvaP3LwocPYzYP
cx30Y6Q9DAQKhZ9i9xrJ3Payg6P8SZGDHIPRu5ZuQWuWtULavO5yfakcoXG4GFIBitCX4mMAcFiM
xleRSpthl1FrcTTy/PIqYyKoJpgvpDzybVarp+v8AgQe9CzQB3AR59HfIKhGtsGedw5A2+sNvASw
V290EbteGqKgsbxjhXJ2tU0ArTgGUQgQ5vecyehOad1ZlTyl0V7wZUPFztmQpXLGCbIwGxoNZkU3
5wXdaO1od7lv3CosaCpPOxW09EbMnWCS5XUrKTtWEWdOLqPGml60VYUwbeJ9ctMFkroZwWZz/uoO
ZSSqVQ6dnK5t84cSE+Yq/TOdznEPG9fZakbSliPxbbkyGowPpG6YJhyTENxsmYmXtdvfLFCZcNae
IkliU+c9x3RaIwzLSWEkf8GvJvLMPFbRjflp89A2zZzcxwAH44u6e2CeMBRFa4Kpv0qVS90JttmC
pWa/91v51664WfYsw3MX2SYYFTpmdt1/GRo9VHJFa7lsz30Er4TJqhlc3FzujMJl1OO90AYduaCM
wt8JeR0+QHmsOKyGLvResQfp++EQHYhntQNs5s7356C+sMe7sWXUN+7pd9LQgj120IYdnZ+EvBov
jhUHjDWSu3DrdN2riLb2hSlyPSds/1lPbA4iUIBbSloxZzu+HiBQjmXjvMdWekJ3Ziyms4GyXiFa
7HHNIGTc2HLbEOZHaCmyCLF6Mtvbf8xmw0RcW35QC7pbt+vx5hJrY9VqZGrRosMxhRkD0IkwPqcx
+3aFA8z2HOX4+AalgOsa0QYkIDfDwFtckVTh2Z8Ccoys9WF3lg6FpzLF+582+Wjw/2SkK4U3m59z
RILI+7tFCFHsmw3WQ8rfZ3gShnIhF3juj6n8hsOUW/G4cO1PnL4qC6IXMDMhGd1Q875o1yx+cEVs
qTGtgsq2qTBH2RfGS9tjAeAeVsNMHe2nMUA0LRTA8XUlU0lv2HV1h9PzdDYHkmLZ8/Z8YEOdP4jc
l8WF1Gy9zUbnZffQGTCT7a0khLofqD+f50nKgeNam/rAP2GV98jsYhZAGMQSQO/vCSe1u6IyaQvU
fU7Vs1PnKbNKOiNOpNjgZfiFOZbEKYdZkwzHonBKSUub4z1PzxXuRXzjO6a9sxUfu2ac7BeIrMs4
JUrQUYfAVZ3/MOpvMrPKknwXwMZRhfFWOpN35rQYyeJgJlgcJGpmtUw9x3M6TkO+bZHND1t4jtyC
36CWi8ZjXDWV4GWNVgCayw/j7ax3hjs1gZoXJhj/mRQOp2Pg9Q2EpH0WSGGqDmfz9aUnTJUivBav
d31upA/n0U+bi9aqOSrkk29jo+0jZZ9lx/32NIC8O/jw2THY1qOSKWO2h5FWnm93sFOax74vjh4N
/Eicw/S4oeIC9i5ikRVA2TfHqv51JMRVSvIPRr2iZrcNWI4tU6yYidta6f6TEPRF3U+CULdtJFET
kmVL1wK/naO3Vvgr3jrmeBBpVAWzkjjNKdli2Uu1Yp9+iBkJMwoVD/Xp8Wevj3m+yH5kCimA6j9C
SkbrOyI0jhWETzuEpZx0isTE2D/QVCojwX2WcVLERi+LUZNxT3B9CQY/yfVE4p5ObGg4d7HT/Ns8
P89N8xbkypIyqr3G0SBdAXmwe6vR3TGuMCCqrBJjnnqMzEw+mBCXD4LKpJJ77tzFliWzxJ+8STtP
jfpveinLrOBElGhzzH7/mm3eFrtTvE4Xk66XGa2XmpInTN+JxAm/dJCCIKijxIBwxbPRXRW7H6jf
6M2dkz5VTtkaDNBuXyPUCkoE0JB1h6/lpZfS9kbdSN5RGJXce2W6GogNzWJbpeDeYz2vbkqM0ttb
1tISh+Q8eF91NtT4f4sg+MB4IjdtNIj9WN6GU2m1nRcI8VnTtDmCxjSN9uxarGAyvZZcCCC69SEY
J+avHjZzkc3h8h4sBjWI0MUNHEqUtc8v3b364ldLxzYD22+FlilslnzMIT9BCL0ez+tyZdaCGMgK
Lz8c2IygzHbwk+eTKWSAXWZOMv0GylP4WlGodhw3WoOIhnHXrxk+WQBDJ3Iif9G44JkCLvTHcEd9
ZDv2iT/FcwsYsNi17L28FexCwcXwwVUs2wuGEw6C9NNfJvjZmlHcHRsKZxaQYIV2SQc1U3V9vLZr
QVa/pKycCLKlBrLCJOl5/b0BAvudl5ijjVnhIyIKrz8QSenEWH0guoUeXnZTnJtAfvCdbz6CgAI6
dfY3a6Ouv1LnqLDBVFFRQsox5kzLsbz2sn2ZEV9lxr4wI2rL28qklAh2yMZl5xiHukjiEDqATkCB
9qiGr4HAv6dULPnO9e39M5rFpFgESdK7KF4j4tcHbq9PxD3x8GYLjeNwNyXaKwKJqGHdv3T2dYv2
GANFUSCV8j3fQoPE56BtMbMgaiMJSU2tHA2VOsdTlf4pcgVCbXTRFt+wF6WFkCizg9EpC5/QxgQc
PzaUPCQgCYtBnr8TNjDnyOAkZ3oVOxLo6KX1brspSWzovEHOE90jBjmELO73fpwkE54yUyuT1Dg2
pRPjDh6iCcdnobSxh4MtieXV9YkU3v8nI42IS+D6sWDVYcH6bwwAGL7CKm0zXhi37BuXGrqsHRw9
Q2yDR2AL3mOibiQ+ZBvp+wFS0qkHyZf+3w9WHye4k6g8c5fD/bHQTw5VWP2zTWBw/9+WG3iZfB8x
F7HH5GHbILuoCOmAVgD724UkHm/41R5CR+JQ4SYw2LfiOdvpz1u+rDNU/tEhxJN930lZFSqcrUZJ
RxL+IP0VcEiLF0Hkl80dQoxS/fL46WgGUH/Kx2GWFfWbQEto1YYovkvQ3AhPbSd2ycPbvJ0lCOQq
MmLw4jscUv6ZY+jf/raV53Dpy+0YUGoHJ+VHHf1dyMMREM1yPMcXaai8jwPtZrgBc/GBtV/qRefM
indIe6to1S/I7TWQq0GI2DrZaOHFPsGvthvAzIC1Uu7v62cHu03anrcaMp5hGz0T42wZ/gWDJY4h
fTCMJOj332qYq7gQUmpspF7lGJqkEeFiyKbpnvwDG7xj8Hv5AVuVQ0Gc2MvWnBEhrNhbBhJQGmUZ
nAqGVNidUoPgl+f+dh9o0tfDAxaG+fxQ6B98aSsT1QHjORggmr/YS9DmnldIgLzAlZOzGPJeNJw/
BQSgVpx2lVlLnUAbtY+RYqqBqZhGF4YTCyTAQ0Btg+qQT7ZayJg7Z/9WZrR/Ui3Z0Z8eNBL7BxRo
czksDnUQZwVQdxL19OYF5ih0aURjL2bKIMnvKcki5G6mSAOJNnLFBrmOc29iGNTiU/bu1mHLvglS
OvAiuH8SmzjXPh+Ur2GWuUhpm9GP5nYXd5tPcTnrdd5YM5TausaUkax0ySgNV7AUjZM5XZv40mtD
DgVFxPkI/hHGUEttM6raGDgAYev9NpwI2xCIguAXAMOUNWC0JiEP8ExtWBqVD8r35vjGTs1S6Fp/
n5kP3oeyjWhI0wIdS4l2cdcgOmplBUp4Vxt0WyahIieEnOfKBl7dac6ZGvvj7DD/1RmivoF2rtab
R04Yn9+F9rpsGaiOtxra1/KabBDuG4j9WrTGjLufeEBh9wyg03LEW2zd0fuJRnUTNhuGEMjGxZGY
hdPRLkURc8l1sNZdrpcem/R80jLcIpxm2b8TMlSilkCCa4ksgI4j6odCt+mf482MiYsaDj186c+N
rxW4i5myQ7LSqmBsmiuPpp1RpHT4hfylHJDgPBFhnPvsJIx1Y1U0sLNRgUITXC/DwwrqIowCDlUQ
cixi18EIQIqnT+ndHUptY7gN1wW+Rjbl721iW+PoA+5gqv84aw/nPDNyH4IBuCOeqvJdBYd+X9Kl
9iU8uxn4zeFX0bpeRc0P6OBlSMd8OSEtSkeabtARToLFrVyhyODv8SIbftQOgvLYnS783kaiXbeI
RXjEjBpbp7bKpz+SX/Prp1+4zeWQSRV69MGceaoC5lndU52hyt3J9Ed0Aki/Ru4K2lL+/6tX32eU
zRtIP+udEEVdciRriOU2wk4pxj5tBrvt/F3q3UtX9ugUn3tUoMLDN8Hy/51oMlQ+4M4/WNEn7tU+
sSpTnsX/iITV+rRLyfFRQmkiclmwI0cWXcs8iFBrf/vdo1n/atU7W9G0uyKmqs00UcD4cnVSImUZ
tARi9D8i4BchJtt9YbEhAloVs5SMMatggwrcVr2eoOwMo0aIkLLmxHP891qYpdyLaUXGAE/mWmuq
ac+fa9bkjUijUasVg0hDMJuvYkTtqgYo2Nat9OIe0VOfUsXes4ExwMlWyHbyZDSTab5KGKD3ptx/
Mog1/Cagx8tm36hWooGMD3SI7x1f0mujXzwAuIUMfi74Ey3jFIsXpmzjtsXMzp0fVcgG5eRGC5nI
nYgI7WudO5h1sp3jRSzB9dCc/tb8n+pZ/8fpetKsbzFJrBBKwA0XeVF9Q50IIUSXRjtJojShh0rC
H9/pwDbk5jsHEypeeJYdJmY26SZeKkU+3/TqsZuTDNQXfXxXTuH5BMiUy3ENV3oBYlu9lTHcqunG
ztOjjSTtHO65oNmqeVJkvH55/Yyqx/vl+7g3+5ZCkcrnCAyf95PGgF/zGEAd34F5Hksb9s0nUL3h
/wSdrMfUz5UVsaX6E7jol+ZYy5dAlzgomKkVByqe4S8wo+LCgwIycDrCn3bJkyI1a9xC2A1zL5+I
MwOMUzYZCLFqkC3T9f9095d2ZAhvJehxKAeYEMfBBq6aa283msxXJ78otcpZwcy7rO2j2i/ghIGp
3/diiMy3OwKNdtSiSdXC/3319Hd0kadGKkwSCnjyJO0ksv1FzNtoTgPYcle7lR1MM+KsTiOOYQLF
sKOt4vfOgLmvAi21V96/p/FdB1GPuuHoWLlsmTT7KSKE3Z9SRt0duChflCeswCYn77i9cabnlSgs
Gx6pNXG45e15uBuQwHqZQpna9NDNg2ml479en0i7ipoAG4upLgcLUrGiosXYJ5ZHR4RYHlYjkMwt
hkC8BczBzmP4s03FU01335L8i/22YQVokcPJc/k1tRZjDO9MVRfI7WaPp5lQXZiJ05JH/cv5G+Oe
DPztLU6PadhN91KWNfPMGQ+c5VDUDkNjYBg287JL6ahjqilAFaABQit9dkBfbIxpd2tKiP3r37QG
xBK7aP8U/nCf3wUAZZUM139SdOKWHrz4ritgjmAphjffIJvd1yVdjFvnONTaw/S/rjAlez4SIyIy
wqa31yz16ckPhYYXEFIc4GcjIYIFyudzEbq9lnz0kn62FfTh/NzPaJ2M/70ElwRF0NQxNWGtScXt
JUBraR/ZirowwDjuqIJfQIAOaBZlSl11xiLygjgLfpj9t7fKNk0Cpvq+BC5O8gbatZ9fAvhEBnQW
8J2X3jQGHtdlY30abDFhXEuKQ54da5lZAk893FasrLNB0I22KCakZBWD3DtvpC8W/5tPsfQV5yrk
xnmDVEiuzK3Pn6qqDEprXGKYiAQPwX9v9va47XF622Z4wsHSFlXcyQ2O8oczRnipLcQ3whOgsdI3
cJdllnsN7Lw+4mm1tt1KAlDeVmDIaLT3HIqJDDe8jvIjPH5aIjiESK66a7zkw9bJml65vy2VD5L9
tuojzP1Il+5pK/nXfsljYa8ErbojwpdP4V5zC+2dmhzojKa2XU1D62AXpEONDWrZsSMVGYLsAFQO
CkknYicS7YQg/VKyKKLvmLz090OY7NSUUxHOZMqL45IMc3n3t4IcPFXuM8TmOjU2kLi+2kXhnipX
q6b6k9aTV+6uvEpNRg6/Z46P910tKObKU/Z+I99UeyvoTG8Ilg0sV7Yklbe31PxVT/b1SdSk8cB8
pzBLulOsajPDmRvfFuIiygpZbBh/tbO9XtOH8cOUXwhV7BDN/85E2ryKEk8KeV1QUypRH4JwTXv1
llRi+8rEAlH6e8+s3N87Qyr3bXBSNrWm6UnHO5gwtDyR84WpEiaLjXTGX9v37gJpjSQd7uWrm8gl
mzsiWrxNAx1LF4Sr5hfzFK17rh+3NCisC6xG6Mrb/CrIU+M+huJrnUlnjlPn/DxCo7EfVjjrq7s4
Iqyhy69rEciw9JeqLtCTAip1+cFA3wF2Po1a1gWgW72zFWLCX7S5oBgTZ2PrUYqr008RimaiGNpo
bQdVuQ6egP3TYAunaugSLltXo6FmR4MWQ0Q77WuWhQ95UxR2YEvph+zkf3H8DljSDN+ZSoMHKFAK
ZQFLCamumY48a7AQ+luD2ItpWY6qbJecoXxrzCXTz5xNBoA2qdvtFUrRrISEs9/D9tpKmJQkSxhZ
WXD/NK/V14d/9zqH2wU5SIUjW/gsIUYhMinCu3rNq8JaAA==
`pragma protect end_protected
