`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UscPXmq6sV0ldGnKnnCAbOJ/OX1VfL5aGb7IKOViidtaNYimBFhSi5UeWnoWf1He
0sgx63YmmwpIeYNWOxOhgctzcp0318lJdPlPFOqD0hJaGF/BR1r5ashS6Jq4F7Xy
Omd3C1adtgU8M37u6avtJ0DPS6HqtgMxEVX4cNIqMrU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11984)
cAMJ2tvv8y6hvMrcDVhmpIoYBRzBHSi35IvW+oe+xFuz8246YhsScaSbvHWwng2q
EDs4Radjti20LEUk1Hx0C0gIz0xCqhDekXKT3o7KvN6WwVAmHZLHJeve2GXYa3e2
Fn31QxmAn5WsYL/VWRSbQpZjVIsohbuYFcOzwSZpZcf87amYDaXlS2i/Z6mspdVC
+ex/DjJE1LFeka5mtWc/93P21Zu5LyLQhgifYZNURbGwhbyhTzR/83VHgGaJK40M
U7M6h07XciInhDUtc3qO9SpSn1EulABxIQQrGmvPo9tMK+Rffqb+3Gt3ryQ+1idr
fZq2Y9QlvYQEZA05kSHg1YBksrMW123MUtkjZD8mZFD4KS1zE9QiyawCGhfOh8MG
Oh2Oq/eF6kN19U/WGbv/43wMw9haY2INy0Untn/4EOdlGDyqyas1CAAS8xH0oCXZ
SebTX7nJSLg7prpxX7vh6uwDcN+37TROLxWmgllp/ZlqDqYWJmcZ+i4STLSPNDVZ
PQPgWJohAQqT82ooVwsJBzbMGJjv89N8p3+fmCQGkGE34l4m45lhBfsPpIDgUfbH
s4HcDdUgYNYsTFNSRV5qS9ONvpJkxqKJZ/wZo6fm+Vu4fv11yxGlYOQZvlk3kwhH
4IwXZT/UvQLhk2aRF5Qx9f92FVirZ+SMx1+dYEZ0Hr5FMj3xlP5+fS9wjnZ/ihbZ
7hxV0WeYJ9+rMArD0VKitXr+zRQS1LaJsQdGbChoTih0lEDXyJ1fWuf8V8jtccQM
fQUVOZwGMxBowJNoCd3w1kJkRaX50EM6Hmy8ZMAomLOzuO16oCjmGPn8VWcGsJEj
7qasefmyTTZlXy0HplET10r7hnqDj0gawbFGjGhb1C9CTV5U+TZqRW9gZdoMa6UN
Lk8wzqq5cZJ+ymt7VnR6FNcKwCwdtpJeCLP2aMqjdNYjk9ak4by63bRaLzNSjOvA
KECBsuhMRohKzdqacV1M0vx/B5vyPWeF95FyS1RDyBIpBedgegTyPvwiz+iKCOTK
nzGAeojEBB3Z4lWZluRAbb7Ln0sYiJyTUw77Vf50XRu5xQzmxTST9fVyI9AJoddP
CnUWaLxqc8HZmjXVAuN9nb14C6JZ666jxr7yMgo2ExRVegCA07aE1b2uowVsmb4C
nDaUj5cAeRlBRX8j3A4CobOhw3EKT2LfadtAq8eyw5VaeL28r7pd2QvMUNc43YzL
0mdJznVyNa7j/KA4yr+LVpUskZVoG0wpct4TMkaMDmTGo/Z/bTCxYW6hKjzeDH9C
bCHro0BPHApBvN1wNH9RgaA1cq510MQ4AiD9h6qNQPE2iCyLTrp2kqXAsgBtJNwt
5XROrV5kQD7ZnxFmYw/0Z1Q+Sayk7oI9/POgn5EQ7SA98dX1aIh+bPNxUFf+XVby
UEzMA5ljIuCfy1Gfxpj/1p3O91yGQW/9URCDjvAd0hKtiZ2ryL+U78F9iQjf7E0M
1EFn17PT/11WOVKIC2PjqQkrEDE2OxJIsznXCtAOpN30RP9JE8tUGfbmb1mmf2zl
O9JWC/sTM1AebJLutytIWaHcBHuWO73YfHz/7xIXPJq5+qJ3JIMirtRubDiSI0Dw
EBJHKfPYYADfTF59I1pbJpdz4kv/CkFFZroGmkJla/+dxDE6ftW7Ym53mPcjsfwb
8tz2RNASiiCi9hSogk1e9Jxx+ZkwszKjXX9Lza5s7IHBYfF3P29V6BDp+uorAI7y
KRcMZiYGesHzPdtNLKnJ7EBneJNkrXsGQR5gQdIrY4u5x7gKHRLP8NngDZervKy8
trQT7Llhf9EYU4y/w23c87y5ziHYfIm6DC1ZQquQKfcAPoZfVa5WbsR+K9zWJq03
gL9eTGVI7m+e/ZMgYUMW5ZZz0wvRNGwG2ByquExmbyP0PUwugl+kuwO49EL1ES5s
WeMtuZxOS2mqe7dr+jv2mos+zY1gxc3poJxUv2V+F3wheI8ASoRUcWaFFSMk68Iw
PZ9gSc/53ypWA8CpWjD5RdK2BHrCt3NQlFankglOuv4vZcjQvtPKI0l0NekAqfim
xWRZvsusRGhK/PlqxsVCfR2qoy3dvBN/2V10OzBWf6R88EC4NEAEiavN8+DvAjzx
ZCgv/YnJVMM/ArjTdVCF2MgEFKVCAAo17sxqcUWaqyavnDaYxHzryPCssuccWKvu
ViQdQb4UWa6moXbIiFGalm5bdbw7HpAQJIDa/XjVc50sbLuLDgrxentchdSrz1NW
YvLVYFeelmbFShxtrEtH1ppVjmz1DS8+7iCaWHbvxUkSzkdpbYTlAPmrcW58L/hl
OUmOEBemvdF3cDcqYlmEtG6xiaeJg7f6LCDsF0TUnqSgqFvhu91is6kPxiMH5igg
ooJNFkpjf6ciStUn41Q97kAZAI3XlqkSJR16f+7rkl+GsYuYyLrI2BKcCbY2MiT5
syTgtFbtrE8cMIJtfiH+bek2xfMMVdIT5EcwD4Iv8aA633BI6OmV67eF6hwyKnLm
hD3MFAALvFevRelvp9y2vh/GViVY8p1JrQz0zDWNjz73GEy2vnSTycL6efvV8SbZ
C7hQ/PN4HjRX82LXIIaHL9WETRIC4cuGpvyXMzXX+922DGoCCfr1rU6ks1EvbZPp
bhlaOUJYhJYDAGDHVNq/IZo+zcbRlxyZOPl/UvXdzZncZ9whvw9yujihL6j5fdMP
myoiLwRZAyd7CJ2QStQxDFmBdLAXyjbsx/i1Z7HaA4gps9sQgYz9FDtP3OjfVkUQ
RbYRihdyuZo07eOq9mSvMuKvYOTDJq6ykZPUVItkNxwtK9jvYgjQmDLcTuw9p2bR
thJ0Feo6ED0NnyhYdmoPyytixH4t259ZvX1zt1r/jJg8+MA/UDNoDDrgedRQ2fRo
mEyGDSMYfjLAny18vQ3MnZ7Fy7PHmYthHPTvGNFM5US1uM15l1SZB9ELGLFOr4ly
I+tof+OQDuDFm31o2nLQqKDWgj/Y5/UQmrFUK3YJIEFg2UWUQsP/fSnZvwU0LOcH
fcafWrC2mf8y1urjbX7xn2BilrybNWTKWjZGH9RLAIipiCuvKSJ0tWog6gJEtzqx
OvJYi5Gku1rHTwaiol5lEdU5i48FCvu8Skd+bCrvsF2AF+XM904GnlDXsLX5HnVK
HcG7VsD8NZFx29coGnKSmtxmQS2gYlHtgR3oh3QyfSBAtaKf17q3n7Sh2uEI2aS6
mIN5g0p8mrue35MeLGT2OEP26nXvevHNbiEpjuKeQs6ToKzWhnOvZ0/sGWO9z9M4
BFL6Rj77crRuxrNTGL5KAdyjVjwSzAOkdHRTWC6/Waf2u6IU2QezjP1j0xEb66zv
1fNXnR+/nFhrfSg1o9e/smd4um00vICu/bREBNmezpJXQYU55tjm2nww7oZYFPnw
PRM+OtRiy6tMd5b0Ae00X7rrZcUmLnMBbvTem6YJ4LAxLy+bNQukbza9eOqfchIg
DfR3suRW3XzB5y83vZb/q+wJiTZ/gF5WoTRp+94v30FKk9fVE8oSuXWtRmnI5u9v
mix/D0u4PN3i6W3UHJV7y3GY1GECKn0FixwW6sSCc0/k7i0OMptC8m2/iblZkHBK
6yiuO+lVxt40E9GpgDBmPZ6co3uTpqI6Cp1sN/QmkylWPtKsvgpjsAVn0kIVj1u4
nmjf7KPZOT3LJI9/CX0oTH94QSv04qT/AX3tqhg84vQ5/wspn4xgI7OO3IQeraS/
Kdj0L/2RVJtUlwgLJ/luGa01n7tf2RznLUt4XKOMdl4BsVKtMtezFrZKt9lDwhDm
FnE6eZJ6OCIM1zqnDfZ5APu0gi1qWEEycw+CNEfR3xr9R+Isl0MQRHY1J45uxZaN
a8v4H4TBHKRKv0s5AM6mhdLVITSsymaqWmwzWMy4ttHIOkbUpXtgnCwhb0HD1lw3
eqrutemB0UnJKm1xwsYyidadtJyCL5ECvt1HUkHlF0nPXUW0K2tbVEK2DBLtOcnd
mFMz+8y5S3m2CzqCkPUP+fTP+rvhmRAopha4STdl8wFPKKBS3sN5eySU76+vqawk
Vrqr75nq4SEAYfWkuUJHJDAPGH1WYaTdIq/1uTJj3iiUhGcgI6aP/ysvzq0MMiW0
+6OOX5b9/WNAYPw8+J4ep8nW4zfZzHknpxSiAq0j7eiaMTQlvYLK7LtBlZRmONcH
84YjOBp4cXEW6t0BAEberavMSCDf/eyHfmCcqJHFo4x3zES55AZ5+jtTsbPZjZQp
nxZ/P6dP6xgQq8iX7jKETqSO8R02phFITaGHikL2jQUsnvRzgQFSbxwBbB8er9KP
pRKHxiarRifCNhfrjHt5sQcG6LJualJGaac1C4vhq5thL6fVcIHD9rfvDPf9gvfX
rvhFCc1gh2+Ajzk+t28BVwGXJJBb7ugFc14DDiJOXOxTbvPbAZgwrogvLF+IXMUT
V9CJKpUc/uCMVuWoY9um+Kfa64U9An/Fdggjridkty3xA8c3jegBIJbiSMzpIhK5
mLef4F6Iz5F+0SDmF6AAZG4n/wQN+XjBaqYxIvFyXameNhcPP9UFfl7nStMV0YqP
D6ZdSBRNaTDkT7YYxLEQq4JwV+OLLmv/Wne8IyvZXDAmoRygLE8eoClkQptXMDGz
ovJMZA4mYMJeBu9gHD592D+OiErCAvvmuUSqkAgsIcyJWaGq63xNBGxvxiK71Lqv
+9OE7r/HByWvbeCISCq+hYHpbG7UINqDjYSLfPdBMR4zA6QKjuYgbdaV/dV/z+9N
RcsbZrRLpLsME8exA7QflmNO7LVZp7dHOC3xRajWACEbLxeJuGQcf6KnFluRQGou
sJN/b70l//21iKFa/AJq/jmlYpAjDCln2WRZvEDoMoEbxt5m7du+EPuOmOJE0A/v
YG57+XwGbLDwBwpqtFDPA4diV3xWbMW4+vP4qEh6WsrDFUAigYTgJy6YSjS2qgIj
JVnbisirQIE+4ogbaiiKFOB0qgLRsTrMFUSSaIImK03V7yFc5sfl+1pWfyFfkRsj
h5S/uHLjHI6zmcggCZ7GIqBjYwNfJ7PkKiky7bfMba22olHRbgzyxwukxLmMc3tC
5m8CvVyr9SDg3MJUTr0gmmlczbF3s3hI5NtkkGiyL6OE9BHXpCiKMwiacL8gWVy1
iinp6WT5Lx8tt3LNP2UtuWGeefVziqe7re9oo0TQM9nr2Ys87GVkHozdCFCG6g4G
ZypnemwNsGl1u3GrsFbeO/PUrdXHQHtwln0SpiYmZntDnd9zi6Bp4KYYkEekKHGh
KhPv5xMFd3XAY4jZrne0mZ6gFk+PJfhLJPG7FwIcD2WtjEAxmMfDeY9D6mtjuD1I
ymltlDKbAJWl6as9N5vF0ir3na38Xuq/KNL7bNemced/qFNpwIdmShngmOrcu644
4/X6+qwEXZtL8KFqxxmg7H/LsaWF4qEZS/dMedtXyc3Zt10n38oGEO2O5nRoJlwb
J+3/mt7EE1uEHQDVFgZADm+aN5yT32/HfAwue7ufBc3a7RCxYxofH2N0Ek8/+BbX
b5oeDpZl5+WtfOC61rrr2+/C1Q99OukkF49gynGRkpkYX09fJRRC2pxrZcx9rePD
s8bXYmfW5HbT8vGQDK3cLeAHppnSzF1WwcN1uWbgDfLgwxqzgs2qgaWaDsKQALJQ
owbGVWmA+QtqDAHqAsOfGcOLG+NBGuJ12axfeNMSVRlkQ6q5lBJRdtSzueNXcqNP
lZQCy1E2nGJdyL6OtAOoAmZZgkgsW9hp1WM7h54nKS21KOwcmkU6sM2D/WKNoaWN
ndJx2ksQ1Xa6aaLAXB7sI1rl4IJmk9mmaFNBi1qwkS4uKcWQORVlZhn2g32OVjAn
6QQcPATVIRFOi+wdet6D4cF8GUYfZYuFYYX6uprDcIjWc7QvL6annTFQOUQX/3/9
VOcnUZt5vTfzSxsCB2FA2vRFpl/FpgTMmU+R6S8b2juHJJYEGQhyU4gObNNLuOo0
CxnlbL82fYvbnC93FOdMAyLNNq5cltBrc1eaTR1h6kYQ2p3AvLUaHmG3vI0AWhNq
/odS75EZI1azcCqG+jQu0E8jfFWcNbbywtrYfIrjrP2vB3fOk8iSlYrPCIwRa3Vh
xVrTGetHmzujVFNk1V2sVAIDISVMTiuhUa1hVi9XdvcXktP2bRtIWkx90RMHvIcE
S3698eyLSdsHIjhpC1bZta9T26OJLiiuldcz/AekixE9Rtm1Ey8NQXLwK0p+JOWv
pjFuxWPYloO/EXMRuZUt0tDZtxVTP8vd8s/klySnADy/YqAsxjPKzufsJNsvMJSZ
VwHfic5iD0HTwNgI/XmqqVmiFbOV0hJS1f3fIIscRKCWdVc6KuW9t2oeuyzjSMn+
FNrAj0xeLjP6/qd5a01HU133NpnufFE+Cdjv66qg/L+WFRMk9b2s/X4fF0AclsTA
ZOf+9QcgPn78J9rhFtC10ag4E2+gwjXqs1gyKOlQ/HFnvHJ6+86JyU7NvAsMqJo1
7Ya35J2LuxIw7zAOK+Dj0mpZ7Z9qJUehwLQykgsRT40NWBzYuNxrftXd6mTOOeJv
ly7OjWlAI5mPBuZxLO2mkGo7KBR7f6ZIfNEgc+J3oeZaWGssmrGQHtWf+GRONCy6
dgfZ8RhHxTuTds+F91cTycJBWohbhicaG3tKi5LjHeNYLLyZ6zjPGrk3IxJCBK8B
fP7DPCg6Xg8pPysKUn5mVjSxXs2s+y3PzVPz4pMiqjsAJP5QAm4p8N3pkywDMJ/j
46C5TyO/ad/R0L5g9h1CRGsfeDLAxZm91nrSZRESCtvgXx8hNfrwG7lFOsndNZuB
pxfVTAy4pXSkprVYnzJv6DGzOx/6zRwp753hdFpp61E2hFbIe7I0Mz9S/D5/eudi
nWvP4of/Emdnagtpf0/LksVQma3ZfJGGqve1EVSIFRko7yAE9iqijICkvW4Lodm1
n80DkoHnHjqceFdhpRNH+WwVxuBREWYwM752NiCKBfw79jAg4559TbgX46mjdM+2
jFyC8wlhHD6/DNrgldGXjzP0jfkNIVypjD2I9fNlvsioeHwzAQPRGq9TLwD6luqp
i86CUQUmRzaku1EJGcElFxK7S8eAUU4zUCotT16US5KXYhrrhvp0V9tp6Yd1V6Ru
3NeVTNnvxM7Lbt90dyNrXDh4uiql4H9aYT8w92k/PwMZDObqH9bW4DAAd8jWm2g0
dZ35EwyMLkegjXXm8LrpTyppkXfgfm21/2b0uIK/sJvKFQqEP14KebkZ757drulj
xTS6Vu0vB6GJTKwsIjmqVIv9xuj4GVrnWzP4MttwaKe1oOZhxQWvMlCxCvw6uY3q
jUpkcyq+MX4xPlvtfITrI1A8ZkkmA7SzIiwCVmGiXTCgfXgr3NByey+nveAMl4Ia
/bQ9qKjwL3nEpuhXEAeM8zZGiU8u9R5a52RPBNiDoEqzLBrX9+PB0seQWJTqcgJw
jSrwucYkNuuitR9vlzB5IeNMYc8/nlz9JMvyic0Wr0YbokeJYOzmhON6Dt5gyPYf
ZxuehGgrE3r6+YtHzn/c1bAcq5JhaIWvj79B7Wt+2JbL7KNbg4EERXKiZMGfdgw6
yhuipjJ6L/3KyH0Zd4w4AWZeQyEwIzONWpb/IOGlWXoxSLxKBsXbhATocCdWCZCg
nSO6YU4fKIlIhZLZXICeF0U3Yzn57HXdXugEP4V+KoSS7wdE/4QSlVPHJi3y7JYc
D3ntKyfThEMsFUYZ5wWpJUVPx+L5VxbC2aj1MlURzf9knzZmXXHaSoCNJWDzbuE3
d60FrtzpJ/VcJW/LZzIc37cazMspr+fKRRgM2PwXffPWtjppCaPKr/uGqVEGx+OA
ERiuqkTtfdGGnzupN9TlU2xGBX/UV7MsOpcWA1j7Iy+3AalN1Q5jMsywnY+FqHSh
uwElXY/BGOzG1TS2hOafTUy6EbqpAFYKc6V9j55L6SYxID0fE3a8NFWMpOrv7jUw
kuZWkHWbYLMhB6+U8sxcRNdGQCoslqdj4SNxMGpWhpTgOkaiekpsYmsgeOn0l7So
iFxmiitgRo6tPeP55vbcLBLT61AA9zL/5WLY/RBbR5CYZCIns0glEqS1MkRgyY9l
ZxSPzdutYVJs3ZxYc9XOYgwGo2v/gRwHK7CzWxf9YqUlNXDrMMb+stH0DWjiK9GK
sGxrFQgeKvunszARxYOCP7Wqbe7BPDCV2fH3Ih42ui+VEYUQaIT6eu8ArvEepsII
jSqbyooUcHI8NnGggt8sgLPoOy7mWcKgaxGtGicvNKzkoFRAdne2VNYDXWHjTwvJ
Sdln+p9YyFsaQeNFo6ZpRj5fh9ksmdhgJtFyE0iCziEoj1hVvm7RiqqmACR/OTJi
KeHEaG7ki12gYb8nq3+n9DsPkegQMSm0Ob/d+5fB2nyCSxLaaQjQ6GZGwDAnLvI/
s5SIbyHLawgeqiQgATez/l9DlqFFGmKLwGqoXvXwZqSSj/G814VMbJlJ4XNCMgs5
xmIvRBmiRYWuVuKOatJNggHUX/tOFPSI/Qi+xmq4JgSo2ct7iNFnMv6Mdn5uSSTF
3NwIDwbweIWDA153K56kBX/vpmmc5MVKPlqm5sZ9OEZ71gpb3180+8SCCxNuFvia
U0acdBua1KQ57Xamh06npVzn/nuP7znkb8brC/GVLa7ALPMBuGLFS22N8wXlUo9J
ybgDi4CuVAdmar0NtAz5R/E8Q4lYbIIRWs+9Wd3ZQoIlORjg25ouHwt/aUts33Ak
GTDGl2iyIkM79IUpXORhTJvrotR54FmGE1pzcIgok8u4AefP19ZvVQgg+g9Lvh2+
xGEU0WysQK2IIgf/owKgrGruHx0VRWgtpNnvtJpfFOTD01pxfa3fdeVlmORV0dbE
1+hYdWUcOYjX03TUUDCYVL3krzkt1K4EJlWnp/BU0xfISrFCMWxJtxXCPj7LmMLe
jmQFD9viXU8s1ovsTy+RK3kxMAjKRZlaUnXoXliRF12t07XPbpT2IBT8QuwDABe2
TW40371LwiaCu9CMYRWpwsPM7nUed4DA+K9AkfFh2yKwHn36Vz7Nr37YWmUDtogA
51w/HHvLzbGw2XuG6CoB2OsVIUo/LoyXKGUd9tl/dDS565aJM+cJVmtlVyq1Q7wa
ksCPqLmt+vN/ZGmnhcAUlrXyGsXfiIxyKjtIVKPO17EvTlM8ZXfnD/2RDyXHDB6j
b0x2nye5EXTa7XNfIi2NWIEQjI7rhczr0883f6gbVnVBi5KxNug32PiD6bJfXl+g
+RhY6lE9PqVLnubaLlt6Vj8Bwc/M3Lx3Ge+6va6tz8WhTCcwpB23B0xAH2vUV+N1
NlCcHbpJJAfNIyVtcSrfwexeAkamvT2fPzqr3IUOQDrzkm7kPlgb1nydcGd89wJv
jVW3GqbmLsRrjiFbhQr3zKgEAuRcaxcviv5vvE3EuwGzRCgHveYxdZb3DMhwqQ5f
oRqft/csVySWxan4VXsKPD/OjATlCVv/JxplRABUzwFRSfsTlCXSi9LxKqYx7rV3
UbuMwkwUqiiopv0CEuhq2lKLQZRr12JaOg9jecDEYfFjkjezk0KJ2EN6twzdBTfq
j192YBOTjg/n8vAaDax0wERdtk6eVaIPyQObmUgRx+Me7SJ3CbvtT/Ef91QoiGOt
WHx3F+bvnQUf4xcY5bA8c0HE/njG0JcFGDP6AMpQ4TbMrcGutKg6O0BF42fvYTyK
BoQ8PNI0uMekmFGNc6oEK55MJczgIt1ocVXPTNcF88vrZtHH3n4fWWm6LijXU+Pd
YZWvXWCc5nxwzZxTr3uZ/c7nyGAnnEBCtej/0xXDS9gA/YJ+qff6O29pM4mrI9jQ
ZKNENH0V18KDgMqtRPkIoDB11XSY0AkEDBIK5t/hx5fz0eVxA3IEq/0yE3oa334v
Iyy90WFmgSvsEw/nvH4uyYs03J5IhMsYgspU1XDYClWU2tGD9N4ouRFPMOeWKlm8
7glBVbQ28Vte9/5tEYPxlDv8ACtPmeDJxJ6YEKF5O9R7QttjeNvu6uhA40tUKtj2
6iA0H0/c9/DDBcZYMnDNG8gqNDZamZ8IEdYqY7yUDIia2PfYTO4gDtiladvrGsYs
wzl4NLaX9bbjlE+vyqSRtjmHd8KLiBtJ5fox0TV1+CwwSfRgzJjhStoTkIlbD9tX
wDn29K07yTNtPeHDZC+g4v7S9lcdIHiVb5/4Aq+/PfT5ho6FUJYI6xf5TGfNCy4J
Om2zjCBEBRloFUW7S6P3X7CUJlT7sH5BJkKn3uXJULTF6StbQVjcSWeZnU5U4SKI
1cY8bZu0Ygo+7QWg+qCJRwaV0a+YVMJeufd1fF5G0jj/H63vcyuhlqBdY32P/Tl2
CyfJ6C1nhhFfHwNt6/iCtrFOGYIreTBwIYsU6KYJoUpqRbpLbVfjyHu5yGR+M1P1
2rxNH0Z3qrUODHkliamBsqn+kJWjZhCTzjdHaSaK4YmZ6LtlSsu3M6Aeoht/75Z8
VrYo1uy0YBSy2OxTF++AHC+LH7TOxsxTYQdg/57XfFOEvldvwoqvPwf2/F7PM87Y
lw9XPGjgHRy1hop4cgPe93EKQk9dsnSQlJXApNU0wZFn3LEqKOK8D5rQTF9LGW3v
+lTp3qrOMmPgwtZFSM8dXsWzWTQcdpEAOf4P6W/DX573H7dCn79Xcw/odnJVFUlC
8cRoczn7qaNKaSYUryWFDCIrNavIseZOogq8c9+CzPrKPTKk7mLPJASugR57fx+G
/1JZacTxDdxIf3goG/uae/C19mcG3yu3LpGumCrFAGVV2nWYk8EaGUsQrpcTV9Cc
PGeu87ik6U59q4In2WkMJYAZ2VvAt1hP8r92p1hctgevxwzjkZyOjLYGcPOaCgo+
ndval6f8igTQW/GDIAS8lN2Z+1/ggw2lxRLWPDGoRgVoNTov7BpPQ/I6hNQ+bTmj
ktTFlTV0OqVQEl6VeoJ0voxL7Rfqok49h/WYDgMgKj0mmOwJwvUCxGIBqIUP0IIo
DYD7mDCiB+zN61x0BUMrbIuq9YmhIlwpRv5fzdDlaJyBctrinOU4burhng/gQH2p
d/pDmBQZceXpWUf5KuM/G1Og8leXQHYEABIn4A4jufWDTggRIIZHhXe1WqQZytU2
A51HPfmKZS55PUQzAaaj1HNTDNiKiphTMe9hKesBmsvDRibtBIA/fQO1GHp31eET
orJMb82btIqXVu9kSBzr0ETUtLH5jeWfANVdMCQEJmwR8he+SNQIqRWqkXEBx8I3
9I6WTEhaLtHMISrRxrU4F7d/VKWz03IvKNWrdlMyplIFVOwYQtLIdHxPlZJrLgPs
XMVN5qAhi1h/BjRRSloPyUAyMCLndvtX5PzecitFzKqZchl1JGw744CjiCqt6AGA
ycCcwn4OA+xBZj6IVTu65ByINe+xoJHe6+JbxWcFbenjjp+xqhsLik14M9gbNCP+
7SDm+bbThWo5QCBe365UAroKEZcxfikAPTYjpXHtXlLgfAAV9mJrNvKRDXdfZxRi
C88BpAgS/Q+0oMnNJ121xcOkSaG/UcU2OoOes/Yk0xZdvkP3LQ1Q3ScvqMWDpWwP
p8CO8bBvkXRY1yo3P+IkYOaWu39Dbcn0dXZPY0U6DWKKjRrAAwMceBf5P6sqpFlS
7jyu1S9eB3rrkjwgM84MAefW52J/MpKPMmEbqhYlxOpu3hkrkUkRYd0cLWY2HE35
m1TcFxfxRzeYyyEnLIHORpAPlpxPQkEEvW9Kt3wWq2mVrBhmiRR6RXuhECyUwV8Q
aphzwI0NF6mS+by+niFrKJL1HU6/qlC87EFdtECKJGsmVPM+X5zdVNB55YQ0ur0/
rID1MyKQiR6lkD/VNlZbU9XuJH8SnbKMOndmmFv0cmTk9LtwZ1+lAhVKbf2TNljp
rCF0KOiIXzKzGG9kktC5lxswmm6qoA/3uL+F1sJzqgn3tPOuAiEdCs6iir/PJF+l
EXsfH2G7Tu8O4ukKJvostL+GHt0LPZDSljWXe06yj9EQdZoGJnqc1s1lxSPVForr
nyYnrXGuJBPLU/CVL0UW4ncj1SP10EwjLArE5BLGEXhuuEOr2VAbxyOb4aspbgfy
UwDWqTsSlVUYLD7C9uGZ4uftVv67ywItfIdjelQ3RwoLyXmwMNwTXkvPvnOZzkqa
K4PjM5dPXX8d2UE6TLBEDjgPsE0EUrZeWlN6MU6A8pfaPV0v3gwF76J8qCG4a7Ez
bgswA4rulMxW1K3ul3mQ+T0Oc/nKpeW5JKhMqEyTaWBQJnk56w21UYAps/oKn6St
gDlJCTRQP0LgrWYLjgrZQDbtIPmtwExhpcfl8S0JvIr43zpRW5YsUEexXXIbw6qi
fxocQzSHqr8OVmqH7Ay+fd/ya66XBIS/rk76Z5L9k4lSgAEhj/7akBLFeh9GE6OM
YuYwd2PIJwpLy9HQjnZV4WZ7JfK+icqInlZ8gSkU7seqcKLVmTOCRrcHEBkLlrhj
uLoVOuY78oaehUGgl52mKCvPBVOPb7E75Qr4+gj/TZ05ieqEErdFI5laeokF6bgo
QB5tu283sTGCyZmM5sPg06AnI1ejh8DRY4FJnabvQFUfYcQglmWon6UxnOYAvcwJ
2nLZZiSWUj9z/TnYfhaWrw6ZIof/BjAP/tv2aNcTmTCJpl/YeSey59GvyEhWdr8Q
Z2GXDLZglXY8mxGINCN6KFcpNejaSmJpXFoxBa1zYLTCwFpRTSgErHLSTyy1z0Ij
rKjmkD+q2PX7nXdNyeN3OwxMwJQFDZIlJMqVv4WARgBxNLGu9yGiHoLBOI+8rTJC
4sXijCWG5pOMBQjKKirIuBn47ZqkAjJPRIC6q+RSYg+fl6BzTsu/KkVPF0F2RFuP
v9fIkw0akj7gXIfMRX+xVJorPaBJL2ZGPYV2LLP9JguJvEcFfu9EWdVfj6XDvrKf
UVfxwEPvK7gVFlfmkCfkbRzbc2J4c9CyyEbnYMS37uc64hKFQJb787eFQjMh8/bP
eZJgcn79AImKeqwQO/chBztTuM9yfkwAZU4G1gTw7Jyua99qKAzyO33SPEZLOpYR
evF+7VGFwakyQ2sEqgw4B72FEfGapy5j2q8sjsKMF65nJMFw/eYY6kRPSKo2wp00
MCFNRGYYYwMV+qHv1vapUpnsEl9ybDVkNTJ6nuhchiUCUbbfzv6PZEpLByyIEdqX
nW5ue1BehTCndlYoOmamdH72MrQbF+KNTbPp30/w4KAagm+pfVqNbquqTEG3EhHV
jGOn5ZEvzc49jbWiIdxyY3mcUVTuzWQPzktcDT7HUplWjQDC8BMVza3EWxU9MWVn
cbyKn7FsXbX+QpRCsWz43Zlq8ijmqGEBna3ZCcTmSeOlpj4egxxr6ThIkJ0Jj/9o
aUKZo8zF75QUQe81BdL4CExiFdwvfyvjKywH7SBT82OXBtpwUiuKhOLNf1VWG0RY
voOG71u/xg6KDb5vkLR04CNopCzwoWOVGWLMTpa4NPaQLqjMpwkpbEinVSo2UQvH
tIc1xJYUJXkThW+Hpq5lteL5IzYVN2eaDSvWnnWb5nfhVFlGGVp4yQXyqVvNKnz7
DtoBfS+wJ5MVNlggC7YEwZIrAhvsMT7Kf2+fMc8+CNisdRKPkUQflGW3GFxHkvAZ
IDXwWqKXTQY6XG2ERAaMpwYfomWayCqSlH7m3otaGH0YKLVFJ5VfbI98NlSEoX7Y
CdR1744o7RLSDNZFpJCBpmfAsZC5XN+aIHIIa08bWGhlqPNfGnY7fXZmm6DpNjRW
yV47nJymMGjkNNn0Z25TVSoKfVogdJBP032wglacDK/1roWek3wDxUObybUdrmUz
MLmt6AoR7QenR+/k9vAcHjmOC/MuuCqxSsbaDxOe2lnRMNX/CECHrqKQJwBiT+Sf
375Zdlm0OwhGsy6ZOZ0UPt8illNlvd3im1loZguaqB9ILBColwlZZlLHCrRbO7ou
VbdcYXyEzs/bGEFmcQLrFepFz0ASLmrbEd1PUhyoF25tzeFlLfS8zW/dwauuXsun
VmGsEZxW90TKyIMg3hZ9Z4sXGfcRA/rC1mX6O7FyM/7uotU7uJFEPsg3JVwW2uGj
ZKcEOa9HDaZvze5feLP4vC6AJT6SA0b9OKb4y6ONDCZphetPa/xqJwzOfFxZPDe4
jsSztIfIJO9uIJ8P2t5l5rsakhCLzpxqqo72iYdAo1RtIK6y1cmWSZ+91htWbJgv
7rsAQwySKmZ5O8S+6KnDVnQ6/YT3jl4PIxBNP4gdCTrCg0LzDhKPsS9QXNDjQ5oj
jNf7BsJ9HEG2uG9iFjYqCh1z6AoI+HjKu4pn9J76rMuGIY1uqefifYeyObBdqUd3
8HuiqBBKxMXwClZDdW8piDJH5Naz1/e4YFDL0btOVlsh8r6gCZJVNA9yVsyaScvA
SAdVqKkdHUeyBd346U1uVFzTP9D5pxmMgFoHY+FSl7/6kKPM4LHOO3cxjUvpKnhs
k7xQn+7f7B3oC41/7+dd2xdsV2XHZY00eFmS7OtvBxReUq0Fq+zc5bfQIAH3eh0r
XWYMiLeoe+trpJzjDza7ZO8manW3iBGxrnn81y0LGDu420KJC//va+ZzBYVqaL2W
PHRzVsjOUjJrFegHVNWBl/DzZJuIBNqCG46ixb0bIhV6Z74z5QKM4SlKA2RNhIe+
/+XMSFkEkI9ExDAtjnROD3Qfj3AskerOmkaQ1/SCs8K1qX2kqlTamh3rXRUauDdk
pVwVGQbP4/yxma4VluC0zyUwQR24/bxX77wHvZe5EFhNMM05FmmBlPBHQ5MRNme8
2mN3+bYUjQk89HNbx59kIWmqiD6GN69D3lOLmLqupoN7RBGffiQf5uyDXMRoF6Dj
yfwgoKtRbEycnsikj46VGH/Ef6eBwvUNbBklUcRqBEOMoMVRVg0GwxUP5rxSx3mj
J7isV53WgtrWqDcd9wWGxrgQm4odDhZIEvZRLdqp4ujVC3bY7r/MhW8GEGdX8Ca2
/99aWYU8im9dCwGcnibP67P1BMqRx2lmMxNkcNHKWjnqFYeilvRbx4o8YUrsI6Fy
HJ1mz2sco9ZjLGEyPxRMAZW3l0F/+dqRbo7keJJDQaUj9pXaeIcj0WI+Jao6S0jm
KkotuEry92UBUeu/Nn7XS0vztGOYotE8WOk51A3YsTaqRmXLZT6HT2bKZGwRDkby
S4lcgtniG1ldz9PotmkzWigqE2kSTB6i4iFOJSDE1dyXIEA3LfBSuR0O0V6c3f8C
glox8yJaqcwVJwpsr68F4XDVPrngp+ycKdf4fnxykKAv/jBfPkF+GcC4pM0b9yQc
C6woAVe8aUpj0dr6agmeZ5DGvYKqJ6MQHVJKaiQo1XMJOmQYe16wYuxemdccWkDL
ZcQi8OM5ZE/x9qhEFe/2VYrE+ovIB5l5FMCKy7WZNIqdN444JCBRUG3B6Se92SfP
+3rB2mR352T0p1xaNnB7fAhjfUOeRgwhc6sT2bpHgL5Ktxrp1D+oobC+m/wiB77Q
Yx6h0yVsj1kkRGLhjasfUX0k75sSySWaTocbE6T0UNoAHmymYMoxNtu0VbUXDEfs
BHXZ9LQ/c76XsRwtN1OgOQ0x8kZ7kpBUOXp5v6Fxp6rBRS22eeqLtL7UZomjAsPI
b9D1fQipTQZlkyg+iSEHGvAPePaVCGOYSPvQ0cYHS20MnEqZEeOesBy7jWS3wljp
AFkDZacE9ml7tmoO7qV5t7MqqQpS0BsQnKedpDP+o2DrHhB0jz1+8OV2N6P6jffz
2F2ix8NmlTcygPZdReqQsrxzqmKeeBBW1ZHJpb21sjEDNBECHa2I2FxZ6TjTpVJ9
bUQEsgx/ikVyuXR31efP0E31+2v5tMR4hTJFMY6v07hVYFg0ecBCvAySp4GWqxAI
RK2KPkbdOS3kBEW86GCHz7UY01XTPW1oaCVmifzHzThMo7LOPrLTJ+N4M9xlxJ33
ZOjtwafXWnv8/d7B4mW8VthgBcRhNccHDGKxg8YZmT/MMCnpe745+622kYFNTL7Y
3QMDzkkRuA2h8lsqWfKjbeoOEE9f3xrTRC3jByCjZEc=
`pragma protect end_protected
