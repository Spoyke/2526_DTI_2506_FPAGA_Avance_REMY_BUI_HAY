`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MAnOGw+vCqxf/LzIoA793a9LP05nBwnRhUUckumO+tH9XMtyXn/ZWBejSxEUB5IP
Z0ssUU2gyds3zGUZtycg2L2sABLUFzinTg+yZ+oC/KTEaacnFwewOgQnIY+Bvryf
xloMOD3/3Dc4sp4Td69MZtAglCfgg7UyJ77x1oM6E0U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 69248)
iQL6mboyiPLv0ASlVvMbT+Jho/O//UvwzgOKR7cvLt/tR53VxGtbk4RHH7AzWdmg
1GyBu6mYA+AmUTQNbS2Fe1P1OtGoVnRYPpZxOGiJzU/xsVBigq5mda0Ms4U5hP1T
hVT5fQmV8vGTlLWHH9SNB38wpmS+iyU93dnYs7KaqmQ3CKEyZVDifIntypj0W7OZ
7k4WTyrKfz2R9S4q5tb40coOGRmHp0IwAQLjq6TEhrOGkm4lXkTFYTgbCDXT2u/y
WljHwemmSzEE+YlszrBVA7zWPpSnfAJgJyJo3bU3Nlf5A/FtiH14ucDni/qtyo+M
z/uoXTWom96vToQrIJSHp3St9WqMCUDt4nF0AqGHx3hL3n93tivOVAtq07j4mNVL
gXlBl6Hw2czmtM8HnuIwoHT/VQ8QqbtC4HzWnq1XkBq/MkpzYYL1c7cRgHCJBTgn
HYcr/WMpQWgDXOq691k1KuHpZVAZgfp0TqPhhHWY2fq0HQipIIIYguMCjYUnU1kr
sotvIDiEYyIfJutORjiz0lZbicl3BwNCpSeg4grKG2FAUf0Ut/oO+QKbicbKiZbg
ZcwXfGqRBQpxUlYK3CD5FcR5U7XlWiRt++itosrBQqP//kHIMYghQphDjVWt8xY/
NYLCvLFVXMy1booiC20XSyemnT3/77z1aZgKweFGxahus8YP7fKIW7McrGaCQj1y
SooVSdXHQphAN15wRPKaJ0cvX1e2fNrQI+ioUsmnSxwXluhKL130/rqeelbc/Ou3
Hwa601cIWGpfYaohIqwoUtBHftUEaP4qq3CeGWF28n3x+cRjepOuZx6qGp9EfVeb
2of1UCVqR+jO0QsKNYEtdcR06lOyUp6IeLjZlwiYyvlaed9STmSM4PG4ybymtgsD
PoozYw1Yz8v2wMB0N+K0fmUuz9x2VNWauI5FqOqlEUsH1ibUS7JJmC+kohnAs29X
wdkSRi8Ht1lToK5Fuy3tGYa5V6CPbOJX28GVFRHCsAHFt8/VrCZ8waAoXgpKZ6Uy
dzVgOyfn17WQHkN+C071r+EIg/yKKY7n1i5njyz+NxL4OjOvE2D2Hbxeiw/8Xcry
8D484xnZcLoMHInC7BmyWQyh0NbVpQ7qAAE7KMtDRWEQFH/JZ8hoGJ0L1olUomP2
ZFK3xa1gg4xeopgE+wOZXDWYByrFsmSTJBq3/gYiPLCEzxjkyENuxgtdbp+h3+Ca
4S3IbmYF1jutQg/z/33i6g7MtdTfXJH2cnk/wi7eoONtfjlXLNg3ENP7F+ZW6dRh
fFizwiuc/sIz1bJL5Sfq8w4/1ICuFuFHptIzogD0ioDNQ7KjN5M1qyu1WZbTpIBG
LYs8v62VqE/+B2YhQfb7QVy9C1HAirn28LEKWwwZNHq9mILEnm+gz4Uv0NHaG30k
M/qcJCcfOvTPZFUw30GRB1vtlK+tO+XlalWgJRs9aEYn2X8sSGHcs+ED5W2kXBbF
BXKLGsEfIpoC3rUV6PXDX4GsAytvNAaxEam1RV7tqBBR7mCpWqmZpKu1lBF26Dnk
7IzkjhWOUKg9u3fyh+6/Xi8qE/jnOZKLVJyPGOQtRwPUKFJUslOHMbzcHN0Khsmb
gbHN+HXp+BRsv10WGMQB5/Pf+F0eqhaOz5KaeYOY8LpuO8U0JUh+8cQ/vFpjk5Hc
ssoBU2IUctX65AfPKzzSABmpVWwxDgkCrbXR0GdKopMwCU6P6b2Iys6xyAC/1ToK
hLmgME4MsaLGYSukxIm4hjNz6PUK5s6trFtDA9SUsViAMn0sRyASUfXLJB+eyIGs
ha9p6XOaXLYNzwz06JNgI0Qy4GfcN/bOzA/sWMQ+W4W6oSYHCZFRY7adGzW/MB7b
D4uN40L3xn5LB4wOW9WfORZJjZtueI/cFddx00mIdbop3Z+0GRT5IDYF/yYHIjTn
gJ/NoMxnPyUC3vQepO+HQiU8ZnQJegkS0V/K+PkX81Wtn4jV/5sM9Gk4x3sRZt1d
c6qws1ZfBZf+mG0QyvKP0Ednh7iECrbsKCN0yC0fwf/mkktrI/0BAaMP+YhkRn7r
vY7h8efQrM2gwnGyK4+/cO+GOCl1Y/nZQ6DkVKj+4d6XlmHWnGaIWGifKeWn1DeA
k3IhbYZkX7S/2e69ZF+VYEYGquntxuisMyG9Y2yOdTNvq31q/6cPK1CXHbHJ8lIt
/lBj0bvkldmqFclEcyYRa/f0iovE0xJdUyPmPdeoZUSCfsp6lZP0uAIXu/JwWblU
OTlzU5bd/bKmlR7k/9vHYKxGCSOfTFBG3FczJpXQ9s5XXvxcChOognoL7XcniyzK
dPUGPEk2fdj32hJunRT3U0gmnAcuuJDWPOVufgn0n7H78fijCSA7+ASLRyg3CQA7
bn2ArrCh4rS1ePe2iO+8rTLFAnO9w6dWfpifLt2rO1/bL1Gl3BkUhAYOB0qSyvgR
t3XIly760OQlB3JS431InnzNKPi221uudBP3mYZosFvzleoS+eq8SYnOo91p617q
WsR8h7UZjbQftZESZu3KMSGCmSg6jzwn9C+gKo14NBq+Ddbl9JZ5M6ErmCmxHcgH
zumc2WwgLD8e6pdcXGqbMI3CQj3OXHPYOMWi4CcExceUk3iiMuCm5MW3TW+yDm4a
eA2PuBAhqnRglAzCG3v6AvMfmDXkTG2Zpi9EehY8QP7TcJP4YL/MBCz1jlOJfv9n
X9HHryRJ+FMa+OYjDawKaUqgTjWyZjM6t9X8EjE86VNCnlo1fGUdDtnWYisRm/Rq
BqdeMOjW5roZE5D38fB49WWjVZMLPA+6/b97h/ljmRIiw8LVRurcn023O8C5eRme
4m3W7qTGso2kELTsMczabMr/c/TFZKcu79biDYkq3LT+WqO2ZNHEGumruqXiLk6R
DDGEjvkEEj0cDQNtONNmtmWTay4qKlq6V1zNbNVNe2kJiZxD1clEN5Xo6UVHMcnp
d75d+piCpPoh418i45UwfG0DpNsPaqe+VE0VbWtCFy2Oufiex3S/b71RPtfi6y5k
46kqIL6zE5kEj/7CHZdceiG+gm5ujcqaK8/lsR3EwhWSMYQBcGMWE1YQ2gE0LAff
hhAASkdDN+y8s8GDKAKbapOSS+bj29jmV2YwKA1JpKaVWAM4AAvn6BqeH0PauU5E
UparO56vQJK+K4z3CycQFhzwrh8fNxeoVb9zx5tKRdfLTY+7xOjpJaM/IOpTM7hM
Qhi31YAPAC2sZQ6ROOqKo2wJgcBAMG8NdIwJXMTf4QePEbUP8gHwNnGYvARmlChQ
LKrxrRtykdX+Xu2qa781mGZYrEl17ok0HdY90gr5lJvHlmowkf3knSond89gukJu
PKkQcRIaPjfaUd4bL+ED1hUw1bjGR2vnWI4PBOqqRcoHO6hDXVmr57QdqV+dvTz/
BlzgAXtkUYey5//8uIwSIJLnGWqsX+Fg7W/e1554lCS9Q3zL8SQjLExI1VUJez81
BMH80lpstVg+hzOTIyhI4gG4bMbPy2Zoj++mzoupsNjzF1T6thJOlwdmrTTg3zIK
ZmwBmGSnVFW8RY28R0A0zIqBcE8hhZGBSt74+23QlCHEGFxS6UIWfLWLNL++sSEk
u5zwKELx9MGEFYXejE2nJJOOuNyeKSsSUkrX4FbmEdxKanNar2wDlaThFK1YYEMw
zbLZgPjeZ5Wwje02kwiBvkdl5DYYIvJOSRs4TxuweNIjxdMd70UPW0mZt5EBY4tA
9r6PPXMIUW1wmGiTLiITq2INGn8K7mBxz98MUi3TXzQKmGPUxdPcBk0PvCpqQ8du
xlDbexgbGsesdxRwA61UBTl21a5tfiJZJro+KygyCnc/dqZSoJlorDv4njSr3E89
zWu/lG0mzElIMMfCh+d2vH4hcAk2bP52tQl1C6f/d/3+mk4Se9iLee+t+9YLOOCx
iLTxX4yq5z+EcpUdca5FIYeMB9ZGTQE1T0J5DPJkBwvM7zzmt+hz6GiujJtOQe0C
MvyERrDLEyEbLRnGIqFyEXKBS/6AkD1ikOcQnaIb/Ep67mp7v4D80PkpamWe5IuB
urACExwLQwAwjgt477KGBkTZc6RxFhJ8poj/skFgPORjVHm1hGoLoLZQsoxQOOfN
9uh0kmajRJhDPWnZCqKhGBLELBg0YDyyPpPvCUVKTVQ8lVGp3jG1bkXfKQSdqaSm
Ua1MPaKIeRt851CeVAWXSnK9KAAM8M/cwUubt8D9i53rZP0CgEVL2z0J8/Us25ZQ
gfzfwqUyAlh1CgNIl4XxJFqCycF/0hYUdiNUIpm7IUmoC1AzbQDUQNhCnO3DVJaG
huki8cpBMlFlB+BoDg60OCnrrqF854zH7ALMuM4I0IZOgK0QLbEkrhKqJmItEtQW
MMieO8CdHDzEfIoCHhixzPU5eK3zA/lZPih8y7LP+GVD0wwL0AUacAa6MD0oC4x/
dkpXpEcoHe6NoqBptY5B/XHjH7TWWr1agcDwjQHI60yyeDe7qNOx4NiJ2hozCflr
Josp2p5JduoAbuGMDlsgWQ+yz1oQT3Da0RG3Ba/8y5ydIVcEUlTxc3eQa4WY8u3G
IBcQcAjpa5N5iKOCmjAigWE/PzmMSUFLMgO0HCWy2/HOwDmod3oK++RqTSmdLFjo
mpkR5rEQdUhWzyHp1sZfOWFH7+SGe0MuR73z9HLq9eJ0ftfegwCJqhnNypY+sztK
qTx9fpK7dUXjilf0ncB/doIrfTB25Q4odFpO81NpqGQM3W4Gv4+UQEVzGOt5eeab
C40vVB5JLQpNahiQVpiDMWzNXDG5TTm0fu09umPnxHjDADKHUUh05gCo994Z8nU3
erDW+m0C/Q65K4uPD3MS00qhNbqOywIjdpTYjMQ9KqmvfKuAfTPTZPNgKqXAlaPa
+9kTZI2eVyjahNf7znK+nnp3ruYNArpUtTo9uhHvSpPAT03X4eeQhBBGMGCoqoih
ejxo1M0OZEgcZ+Z8NIT94PPlIxWxkLkg1Qn6xApfkTFZZ3Q7a6ZO1IAoYmgZXFqB
ycMkPnhAp5O389bZWIMiGR0eGSLcNGBGyMGDxFl+yWatTvRzUq8RJJZOB0gXxiJi
2wYZq9gRBemIofeRv/OrclypVTa5PuJqAx7tCyCh0EaBRsCj2sr90CRDxWMmK8Kf
0K3dUwEBszvP/kJSpdAxjMpxPzQpZpg8Wc1CmKiUbJIKKZ6vkfHFFVLop8g3UOnQ
miwBNzqlm85UxRuWyHBcdzkunscK/9lCLbY6nLHea5bWr+xTRE0Hpn17voa+PDCL
08OOfn70iznNA5R4hQ7y2BUvnGcrijmP+1Fy0JMn/f3qVZRZeBV6Js8HdRvmoHiZ
LgC5D4vSWRX/V1GpNkcYmtXmIZ1ZpHPVxooN3M7jjRAUdX5H11ptqAtsJ/UTe+Ox
9znnzvoQ+jDxHmYiE3HlG/NWqAzi+o2OvFKzaczjVm4DoQm1TFVxQgmJbrRb3L/d
XOncV2STlL4/QgNTClQCPJmBogLq70nIRh8kZRDCubfR4JKNVEaIXuK4tplzoCAP
s72L9ZV1u4USpEjvhvhEtdiQz3nBxs3NdtPEAu1JCcRpBJJIHQCIaUMywakbDM4j
PhY5cdux7gjjvClClGgOr4WOqo2OU4168hcZVFlfX+7IjDeUeaeluxbM5FwoiypL
sqhWEE7H9pipKjiQq6fc27wKcKHmXZj4P2i1R7yzk6bd0nkbXoq04lq2Vr3tOG/a
6evLpz4690+YIOP9BRy3cFqV+l47//WCZeSc260bF3nh9tFrIlM/3wEJk2n38Ub2
FgAPmmSBafMcVKJTA+liI5X+H9iWE4pJy7yz2PEivCegB97iH1Edwnn+wkPR/qwN
SfPq3/hoH7bxsUnFwe1RGQ7R4XMqWUguDzncL3qOPosWLboiY4EHMsJqzln3oDie
sjQ3z5r/UY+ph7lpm4rjJvc6cCFqsMOv0TW19esMPhapBJZUuxj+i+pkyf5Lqi7Z
FgYbFdeC8lW1O0kokTwCxaLznN2Z2wxIqYs4bgpaM+dJEJnS53Vd3gZ2pzlupDR8
A+aGyh3rEN4vVueDo543OTGqAUpHkdrOEmbrYOZI7VStlWXyn4r8sXso/vl52kNh
YEbYZyojvZQzi0lFnPrI8JAEu8JFFCTRj2uY8cE0iIIkS4JtslfnSvppwObDgKi2
MUQM7Tx5DWAJjV/4/jeqR7ZbB5NjRvkK1o4CZXwHgxXeOK3j7D61adEVby+Jlafz
Tmbb1TC9pQRukpACYe2I8ttpwvStBxgiveMSVQYoqz/HgkHJzaZ7PDCrn4YqE5jk
1O9oIvKIZjs0bsZs2gwEsicLkhnQBv7hpynpKZP9OmADzHHOYDZYdMvyF3e3MqSI
3wroG2gGMU77YvrobkHsJ2IaCC2tL4S82nQP2cJ1MG1GrcX6yTH9Q014Khx65v2E
Yt6Nz4uwF+UEibbiFhGoBY0udKhXjFC9RrnFYjTYSzzLTQ4scTz+0Ff6cclFXmy1
d7UrXe3wumu6NzDWX1mYGS4R7b13UP2YxR7COigNTeOYRdhFEFqA5mfYPGMYSw1S
2gF15bTElJKfDk6UvpI49OWUvCr3cnk2mDeUTOMinZX4DvomEe5OulgRb+Mg7TVe
Wd1RGmwcCHPvDYSccXqExd4KJ6H6LDzLhce7b+CxHympWtqdJFkCxLrDGaDC79ld
fcf8yr5flc0AnLLst9p0+OjDpjY3NilxRSZjyCFGcxrshW9bLdpoWE+mmqrDvWrF
rlQfvxX/nlnXaeCkTA6UIiHPOgrNZvFV+exehKIdXYHYbAX7HRDnzfo4tQ1Sgr5q
B1nWi2L6OZ1YMOHxRtwZHQvjhejJs9YgG0DJO5FP/wquEwQHBbWH8PYZiYO+PFEa
zF+IRvycj61EyJ2AQ66HMicMIfKn6AMdAXBlZHEtIK9wsa6YWLLLZbL3juxfFIld
c9e+T0wy38CHDBGm5FuZFxLlfB2BkRt5jZaQqSRo71duJuGhpvY08t412Igm53G5
qDXMGOIMQUM/Q7a9/1wisd6OTyPd0c4STYHhbUKgPljJJcs4h6Z1iL/Ihap1ms7o
2Mhte+BkyIb6QqESjw7WwxoFCw54EPuRCJz/mdE/DxpWnNu/NUPkhdbcs0ZmNLT7
631blhXyMYMptmJhz6WnTbj3IipHx4HRJor1V6g/UB8B+2Fu2+gtwLQYd/6l4pjZ
6O0qQiUQRzCGenlHT5z9W1EAfSVkkUkLSAnVklIIe3CT/4aeoy+iBZB5kBbGtRzQ
vQ2LHY9I9QbUSseaFXBtV86P9kU5wzSkBeiXIsGWXYKOI7XqMTRhBi0wqN97XyW/
mEbgH4R8JQZ9vCgO2geST6MZOOuj4PhHez6NOzBgYyHywRNLNllQWdO/y9s7NAbE
moAvcKgtO9T9ahG8fHYABetkt09m/qFXgpPXamhpKW5JGDyd9p6ScIpNuZas20Nv
h6feM5mNgaAvB0f328OTWO4wvNAxPakIq2v0+Dn6G32MRQv/HhrXFzzDnRsEleHf
mYcQp74EFX5q6s99O1IKAMlG9Omuz95D6dcjVxC6ZosnvyHrewkLDyh+gABQrfjn
uAYY+jQpIRTQrBMc8hVFgII5w7NK1bJvCQyway6zCNugFR3JAQDalt+3bagf/Vbl
UIWdWT/e5QVT07JozNTaACYNqcKoYI7cm4lnUueya4+fZqGDGVMUGScul23GjvFu
1QiuwlM3uthv6NgzE2jE1ronUtS7iCb6tJIcgeCHwaGXXKU9OfCBb/mbq++gShqR
vnb8HS7SVTXlanUakYA1FqszWuPr+ONGQyViw9By0TNlmYZ7kCvHhQH8RsYo3P6b
L63we3GBPI9dOol0vV9p/JlEGD1BFAA7OYRA37WIf2Pcqci3PSqimDh8iW0428+e
pSSE7uT4vzhL4Gdh11GF9nNnIOpAxx9ni7IEqBDHh+bKG43jVyTiPkpZ0YjXowI1
Chb9DuzYDzdBzJMgJ8rfGARNeOEMcj1JY6kPM/2/yPeeVja2AjeZr8xj73rGjqbD
8HDwFyN9Xlr/B9Mo1aFNPOc5YI4TbTTHZoMUeNq+7GOLty9KkfqLpK7ijrtdFa3w
l44gQqmOmhhFeYbRJvPyDQ5tNwQN8xTChGXIpxKT54aCn7ddJjlFVQqyS1mPiWyU
NyvMGyB3OdGHB6NoAcb8BiF/3iQ5M6DJTIts0IqyDtMsR/azTdp6stZ/WZkVHkJY
/9hXXlsa5TLm4YzRs9HqwUH/wJzxVJ7d6pwNdfkTD2ypAGZ84V08V9Hzg+NYWd1i
MjuqOZBc8efO42N/W/yoRMZhKWAB88aMyrulpdMx02qoHfFqHI8zMQypTRgdvDmV
2xn9Hww+goQhgeHAVNyd6vvcKDKq9iND0ZxM/+BfYQQgc0h6YYB4tqI7Rj0lmi9Z
EVjWJQvPuqusYMS6yB3b4q2kp1dVIArRBGbf4P3Fu1FixIZl5y6D3AdbbovI0VvS
1GVtkvnK8E5l+cZwow2gLrATwLDpA+wAB53NjixNO3L4XDd8kwGsmg/HC8weCc8P
qoO6MPR6xl6RWH8yQ3zK86K070M+BDLj+FJl0HpkYVgZRTOQUgNCpkB49nH+62e+
ZSMWw1I3gb2b95IkPy1Y/FEkASxAYgiB7efHaKpy3tqmCzJ8wdP5237sRaPOy6An
KmUFkc+4+4ZoDeB8fHw8+b0IQEB0LDlH3OQsEA5M7Lf+P9cCA0Plr1zAIclNEoeU
sViH2ta8XyIavIkdinpExh7Par83ddUKV/4JIET9+A6DNqPrFRc33cijb0XtyROy
7/gHWJjBkeAneeZOz8EsXE/fokX/sdGlMTpdUFric8b4M7gAQ8E98KtvrA4eAlT4
nsbPklh/GZ5GDLb0RqicOtvFQqj6IXgeYVpvrnYJUtA3ECzqW/ZH3bmtwpABrQZH
i2D4YUDkbX7ciA5en0p04HqfxrPDthy8q3GCe9SgYTAEuGAQG6Tf1Wgh3Ee7tiM6
xsl+0d62sGbspB+jAtW/PIqG5xGDtUwMUfMNrKYbQE0XaEV+JsenZSOCbCW3lRlb
VAtlMx3C3WRdc8vu6eWM2E5gFQebT3L+9Gb1mp2TaLWg4mgcqfRtpWDw2zZ5BjqK
c5Lkq30RkIB9ZoFTdkUtU/tgNz2IlaAxgl98EYwmfvPU72HMHV+RfWlAT/wFo3Vm
se5NcmBZfqJMkFxJf0qUtHg2mqJY2prYBWqAqw6vMsJ4DR2HNYrS5FF+xSsCUVeU
s14NxA/0HgxmvuL/DGdWCXDGmoUfPhqLlF3cUBab7FK5Z8csRAJw68eyGZzDlY4t
mv6X4qd5oUTkn10kPbPNKvH1yojZesjJGUostqdY+8jdoiv+OCHNVcjLjN7rT2d6
4DpPK6K/KL9IP3fRp+/gC3kZqGcfPqgNwfYTLQ9O0U9sV5u+lI0V1GP7SrjdkrHr
iyhIC+JI+2S5k0FwOJ1e1X0yDY84EVIkUkqTeNI2k7dwNOSaZO7eSfJEuME3NeYk
d+ilTeLwVM5BnEPVopgXohKHQmNZcAbMFLfbOC/oCPQ5cJoqmDJL/+/Oj04XOlTz
NhZsMI6VyJ3IclaUZG9vIKlbGrzX3xQZfgAwXEQ2ka/gHUzCwp+dFvvWQT8CFBCV
cW9GLMTBitFbfMYmZ1Pw38Ok2LjDn+BAUlD3b7V3+EPTAlMJl8/gQzVQJUr17ScW
QNL0ORHzsyIkcTf8R+A9TWLK1XiTmE/qv7RpomhEp0eoF6tkMow6I5IiBR1I33Un
EwX5B13Ioq6Twlc7Fal9Tu6YeLRGLgWg7TgHRzbkh8/2Efvl/gTWNUiIw3LysDkB
Tj0+cIvHZYuuJPkg7WmIbjTT5jVvC9iJs0Nl5ndB0koujilX3q1huU31VcmBRQB7
c6pKvTXpa4J2QXNzJhsBL+RaS6kdEhYqTnWHHHMsU54DmcCdGb2I3oN8eQBr/Jhx
SY6oeX+1DpNbt+iCBXt0kUTH/34OJEnrInhSeOtpIReYW2OkCsb2WvDcEYMVbemr
uIzCLU7W/WLp9Oo3VLGKzpa046n7gfKVzGxngmeqoP2iEcBuIAzhDSsLXvqkBpPD
3gCkxf84XBZLYmkNyychCFLvGgVxuUA1zZVzTBSKBgHpeqp9QS0jVUO//GWTcmxc
K9C18ehKGW3Rp0K+Io5juTk9jVrnVCLYDY5dErXTeobk0Gkvh4FtjcySYnHNPZcQ
BE1y1dkimT9dsGos5FV2j7rx3nkQ87BmlSLv0OuuNqdtWUCL5IPR5wK2s/1gufvx
vYGzx+uVXMZEuHQZO2OvZVj4KuyuxTnXMasMBN6z02bFv1JjWD04aFnJUIY1uGIn
mchdyw1w9RtZnnpiJqkI/os49IrcHEjUbah6IFd1Tfld9yaDKAuI6ZkvehUbKm7Y
qZ2wApKYvLBtVXvkaWtm4iSFL6mqyFfX3W12fgvXCQL6TlUWtWuwzSmVjeQMM0Yb
Qov4Ji8JORQW8CKYnLKZt050DgE4T+ynd2ZbFYwh09aqtcAU2kiT4vA2QQ5ZtIo6
8sIMeIzK2AbglRL7ezIUpxoZGfUipaJjB44QYMeins9hdMsWXL9p313BGq+nhj6K
UdhMYATEmVNeYwvdu622kHs3wvyVJ4Sn8aoleroCt/0LV0kzyIDIZKwyKYvTvkQx
FxoAVYQYQOD6Pxo7oidhApaZ5cUWXrCLquNPwRZWT5Fz5hY48x9P+Z7k1tlpisyV
DiZhmLqUZbvukYjuvFeVLDiunFGR0MyxjnGlYwNqhJyMDu3TooIs+wUKbZcMU8QQ
kjY7SQUzXZnebZTEbtndDnRFv2jyUXbX3rAKeR0hZIQY2EnxY5tff6LWfgj3pV5Q
VS7S9DxX7kvX8hxYi2eyqwK7HPbUEv6hF6DRUYsu6tJsZJ591tpyeGVQoDx5d1eK
kNvllhTMMHrTsxA0P89itJm9DL6iKS/Xx4fKaaC7b3mY+A9/H/c9hRdc8mSD/S7A
JgeBFNiEmlywc05crrKsjLPVKyjLEsCUIXqYm0ZbYS0aw37DqDDtwkBzil843uub
0S1edRwdgzC8Y2FFWT6ZCGZO5xYj8yzjlv9E/6SPEe3k2FGZmzKBnodRsyzoVRPO
O8wbzuDZmqBE3eapKyMWMXzHgbFpEuP77AoNHXQ5DEmDp0XtBFQ7xFI+Wsw6ORzx
NNPXV5feAi+YFeY7azUEtcM5sogsBY5yFmAjAqOPrW81mSHpoSIdP2poQBB0+ZXv
wClHtrYN8dXlnrzdK7lCPzlJPcUafQisL0rCipKWdlqMWeUw4Scnk6JrlqQyXHNk
iq83DLrt4dsxfr+1uzzsTqtSZ+1Q3ZDbDtNFmzhxaMLdtoz6jDVYKMoSKxggkxWh
yBRY/ShhfKEwbYfXMpgyNMFlRQMTpp2l6x96e0jLN/mZlMeRe8kX/0a07d3vsh3j
i568Ah9gfGSWYB48k/AqtHyd5NE4zh3X4JRXjSOVVUF4cVO99JRwC/nsRqmGndim
wzwMvaVkYGNuC5jYXssj6GUMsMSFA3ZwIhTJV8aFd0NbRipdFejB0PfPU+rsvpHg
iWg+7djH9W0DEnfx9VBM1NFUthAzFHqsAJtjT7aAmFRpX7uy9uY1kItF8aNw1AdC
zVOLO1aQeGicT0bcat3AXyUMzWOIBSzWdUh6E083xNP6r0gy7dCPhJHH08/16gWO
5ZbG3oh5pggMSLYVk+5lTgifYvXRYdueKFX12sLSlTZ70jFwCCOstW8Jtwpmyp/+
TNVOUSzXLirGvTt+xliI+F060D9RT3YPJnPgin/lU/4P9TalQ1t4vj1C86lM9zLe
hF8xuYgqjxczHum4sJgUuKbBJoQQBGBkXOaCVf3U2wlSk84anmnNWe+KS57ESPJN
fzgd4DuWXN4p3jq186OLfAYPAxuTiTtELHVsXNuql1eiT53M+vIhqxuUoNQOmGos
gKxK6qyFysFR6CmPJUx43BtcXcXjmjnFWkydFu4CgpZcXQMY13TRdGBoCh2qtBxP
peBX7gtd+DVM6+l/SXiwDNK+DERoiUf67benDhFD9banN9D21ih0roW8t9h/59cC
i+Eu/f3CYcRpdhmLP2PUppn9rmN+sVEEalvd2kPdTf5czbaioibJwd8aMUpBpzx9
tr/S9rJAoiMtZV9YQ6f0cv32lBAGZkvM0Q64tmhftCaGw7jpHzJkvX+5KHtwvXyB
TmmbVi50UtG9g46Phzqls9ev0sO8yuMSS3SnN1gJyRvLpITbV6kpJqXemWKC262c
rZknEKTVOXcbreVRDmbDQmZXnuY+7QaDbTvURT1OAAKCY2pY8k2NcZhroxyL+5B0
XnjZzJc4tsvMRarMFDDknkjIzB2d8tCihwmScDwk4HsLGM3YNqLu9HPCGu/HoE6w
z0TVynKlgtnG094DVi0nH+KVazsDpFuc+vN9yp5j2qj+lpp01i93WIIPaFYfYA4j
r/IfNo26eYGCBB7CuNaLMGpCCK/BzsLwl0NubIjgd8r4eZRjivsewlLAYI6of2RI
wUWWLMkcjY5hgZv7q1z4BvGlro+mTY1n5i2/+vNtEMW7mzv+knTE+AVBQaHFN06s
pfDmVI+H7ua7BXoKdkdDBwijlWKa0CjVrQ18FRFT7PUd2zV4yxW4u063hVUGhXmt
QPw1YbXJumsMhr/XSYwm4eo71kODgniT8Yh/aaejRgF17JE13fc4KyLm2duSdd5r
jmanpvLY+sLSiXuGixKhN0uOWHomNYjCTpiGQASuZ4qkUB97TedDb3b5C0RQ6dnv
Fc7nDhRr27r728pkByQhfSMXRvxwh1CMzPa6+rDxVIDMhGDtd29fxyKNr7adab7B
tbUrTL1aRWcjmOOKtMfCQpXzGX4YsmHt8A9dpRYjEVbK8ECUTWI23W640jHv7R4s
3at4FTXLv5YRsoeOPF2qjlXrq1nixr9tE18p//C41o83S+gKh7LZvupPy8Ujkd/2
N1YVpZVDF4wN6w9WrXiVqbiM6bbOt6O8+p79cnaQnPFh3YdaZy8CjUVyDnG9xAFJ
PkXoS1Sti1VN6YSMrE577+JEKwg+gF9FJqwoG1k4FVR9NTtigv5hB3ZvWuLLFBh7
b+6Ct419pfVdNhwFGrKgLj4R+HPH38suV0iKD5+/Qd7/XaAycy2j9EoNufybHR0J
J20YcimwgPkLBV3KT/gI5ekGEkmIzd3GVIVGL7nA/1NF0bIEmh4dRXsg4UOz5KYA
3BLIMi94AwROyiQ8vdcyWNUjjt2l/PYwn5gA3K5faaKSVZ4RbC9/P1E0wKgjlmV+
AGDF2MU2wkIIL8ei+/C88KqRxQECt4k+3QFhn+Z8uI/7ChZUOvGAfTHIarR+cxxG
Hy4rwBnK2KGzfR4OH+PdbM5+eQW594bPuLPjVsf2E+jfAdyWamifU6TQZOnBBLQe
Jcf/ntvQiDU/QFfFBsY/UBh4IFvw9pl9e1QtbIALhQ40UtOeLc3btXz5f2HAv0AS
4byiVMpLTF8uVURfgYUvMYA7h9k8O27FHfq92OaLZDDg52DLEEC89ZEME1RYVhqR
tgrVT0lQjoLT0Cb+VgHRfx9ihdvz/lWOkeuhQIlzXIYVX2g66NAj+N3Bd0wmyvDi
f4vaXepmpNjXA5kxK4zL3HcFld9ZulDqIr9TNlgzgVM76JauqkUxmuxBRofbTijR
eIWzecDc5W4sz4AdvTCQvm0pu7GH9dJktf2RUjmL3Sao1gIlDmhrMgqFgU6yKaSd
YlBjpm9yt3mTR6T+zSr7uYmG2hRSzEQnMHYDw9f0Nv3LOE/YW3uAl2tEPIx6rFJP
l9+narXHOAnKNsdkpmDmJhEa1tF59AT6Cofz0TufPbPFTWnKfGhI6s3NmX7XjZK3
xU/2fodC16912c14AOgF11gyqIF0qkC1npIhhlAazx4E8pXrZzPDVFbjGNgJZmQI
w3r4VQMCJ8oGBele7Wazz/x+fH10RQAMOxDPasw+FiyT+GY8NZ9eAM1zx+Owo0F9
ym73IdvO8DvTCmRKFL0Mg6bLfI/px1eAbLa7mK0Z4PNnT907mRezXz9h5tx7Cmj+
ik1+VYvmyfybQNHaXDp7UFOuaPuKpHKDu6Vq/qmPba1L9QggmJgW6UHQXO6HX1ZN
HESJ1+vKnfAElZ1dNKnL7qa05Xa3AL2gY2y7K9JaduVOOwkauaz7CFsH+03XQwvI
AVYM29Z+ey6lxOmiIta/SA6rwXKMy4RB922gczHq5F3a/L7NGS3Sn2UhUbN2y4y7
8lXlk/2JJz+7d9ggAjhN5Qe/dq2l4vQ6AVcDbl8gkgJb9vOvZ9Gzr0DcwhDRHCIe
OO9wAbRNdctmUJdItUbYVkruOcmiyqxmS14cFz20ciI+Z++MYcz8g0A7DG/jnbLh
3Er76AhFJqw+ONSOCrTs6PHpE/phcZU4GBgOGMPiTF7e9W9wkg6ljgmoQgSVXSDZ
W/nVwA/Ee3wLFjuJAZeeTVIyy7n5xDxMnPE15CN4qPwtugZnUdd7knFUsAWSuXDh
pZ01Ez7EiYOKnkcI4aaZNAAr1Gt2cKq3wYYMfg7LC5f5jaNfZLPOOotGVXwP8vk1
1SN/RFtoY8mQin2zH+Z4W27Lt3vyMSfwq/xum68J9aat7AeM/4STAWtJhRyIBP73
wI2qKv4Gww4H0v0BTc9/pvptlTJjk/yXdQfdaUNf69k5vdbzHKhBpycHUKsEqYko
94M91CnwymmZquePLsLgXlnwRnTjMFApzBNgHHzUOTDdRc3Yw0bDLTrG45PSktaR
7VIOqLb0vZ5JPUNQ0CpToRWWkUqYlDKMBQqfCJoAtSu9Gn6iream3KpFPLVUw1rz
rt+/9+53wANn1zXuS9dTvF1JYX/ATpluimqOlQTnz3ArAJJFaaIw0MAycIVfTdjM
GU9hBBp5VSKMwATkkZJhwR5yY2hKtbl65CQ8p8gmRWHuwO4m833FyX9eQWJH2tli
6+IfucEj9qt0yKHFlUmNz73QXyASzABO34fCw1xw+UkfXz3ND2ZmJ6FbBHQwB6EB
Mi98Qpqp/U5WCG0AsJ4A74pkvzmR7t259fTtEc49ulUe67FdswxFjPpinBFh5V36
J13VXSx8/RmaONEp0rFglMuPZRsERwrLMzbAv1mqZRaEsaa3/A6eMZr/tPoKhFF+
F8yoBYU1JMCv/lPrbXGrUJdXWgmOEkLHc/69/AoyisIcsv7Od9z5XF5Wn7mL61jH
RGUMXaoejBZi9oLbaUJ/Jy7lQR79f7HbtMgv0dti9k9rreZhR8fFlVaFaXRzJLEd
GBbTd4o/ViQAPRc7I1Zjopzxf6BLNakLWBCPs3p7ahB6MxvqKlFCFjnh2SDuo2vi
uMfW4Bv/aJmG31SvP08s3L8mtL80NpsmPGatiBh41Zl4a5oiMLjXPP6sCEVRQNzS
SU9uI/VYNXqNEqcCk+YAGIB9GMPm4iuxL0qefdYP4vOHJ6ByULaADjUxBAgWpNCz
lv8xxK5eyApIVxbeuklI6zgmN5AlTLkLbFjQqg8oHz1uVVdBUYMWUZnBaFEnCLTf
4BGczoMdWUlliQtW/+nfu3YSZ03Mx19DUB/aucNvO8/bUxc4d/Ue8p1fiu4Yt1pN
9A4jMeJJeB3f6LwMRLEqCuVqDPcjbtMRacoaqyteUxaGUAOZrh0DYsHlQUadRZNE
Adpz5pVJy80xw3dk3+oNZqsMwuYo2B1KMjwKOPh5kAnhKeYp91uSnKL0DgbbKaLZ
Xr66S5FjU++W2PwF6rD3tOA91VN+g5+sOHKqLpYDE0ig35eV5qsPx3DehBT77dLV
GiAPxQ8/Gllsddhha/zAyJY722GByZ/L5Qr8cypl0XjU34FwMpKJDdaY2Glfq5CS
hzLp0rl4gctnD/lPY415epcPRPzTjb/ixVFbH1NvLgNUPrhGcLZTiSP/B2ICGML+
eYuHXCQdwxM0AYWhZjNvXxyfQY4TMOOzvgya9TiyDOm6oFkEhIwUNKvZZi0oZ8cR
70AOLNNL3eamr/PF78TOUIrZiP/Hk/jWBGHZ4x0t6QSDenjCY4cj79pOmbcWPivj
uSdTDtF+BNHjzeB2xkj6+t6WjfLDZx71lB5xMivmqi3egSNuQ+tsF2brnr9R26Ie
smNWTLV5cIAwqp+yRSShxJ8WKjNnjCxtYPMxMFfIoF6UC/0dIgWjuju/Az33sX68
08l4h7rUZpECDS99fNdllFq5lkRFtvvyLIjAHcuaiOmABtR2RzqYsbUJBi1NcZz6
1J3kvXQQcpng+j/sV4IQ8EEolfa2e16YDFMuGBFQPamD1ObTQMa6NIlFk3B+Mn++
Ahu+C5yYgx1/p9O6txWwgxuNRfZZqPkv6TM2IQVClGmHRAwvDx/GNRnkY6tgkmap
j5uI32vjvmovwd0wMJsCMoBLZl7IDl2ZaslqSKWCsw4LcXg+YAwc5ntcR1vbrzKa
PwiCPcAIzha0OcpSuoc/9wjAG23jJLDUBTYPynLYG99cTFOAwkJCOX1Ztedjh4zB
3L2eAnwYHye14IgLVK0eDb8dsgAH9hLI58MoZmAc4EWYx6h3DvQ5anQWKpg6jqtK
e1HY2jjLIQseaPrYpxmedjihLxfvXRX5yUBuja03gvYv2oWYGx/M+am2wSjqZGXY
pkpN+P510twECQra9XtqDeZL5XPGDzdy2Z1U76EFwbWY/y4Jd+WcmFuBF20hYyNL
npI1rBqk3UK4v/vuadc+sXxs+VUuoyKCUk5Q3mhpAPofsIcAx7PfycI9MrJ9v6k2
40XjJWQiIv+vXKOUaz3RoG0B46UikqHQP+kwt3cmTzyJsm7UU2VX/fe9tYETrGFu
dtmoCX972xOS2ESOU0WmGUwWlicoULvj3gkvBs6Zf5r91WzYJMpjAw6dUt/kDiXb
EipuJ3ocbxzuyBmEFWadlOgxhMugpgu5oMEaQWOOMRu1j5ZGwtv1S1AFuwAx4j8W
FjQhjpQ0eIV0SOIz+0DkK3Z7yPoCiIgWMY2Gxkn26y94eQ0nnj3PO9YXiIEx6nyH
kom2gjD08Z7qo2RtioH0YgQZrArQz84dNUd/iVk4VpAIQXOLdMFuyHEXjaEsEQwC
XdvMYdzaRTGCvfDV5xffFq/1B/I0PCzActN/UGTFHpjM9ds4gzy/3zxKzSEkBl4B
ujNGKvKx74P1p4BqCZuYC3LqPYE/kk4F0OdhxF++fEY9UyDhzHDqu5hATDSZLV9N
JLy7PjixPc/N6YGWtfV/rdjSsVD0uWlERF+RGTuGfs9g6GoPMpII1F4oe3SJujRU
tKrwEeHZid7ZaHAW/I6bUf7Nm6FKiskLN6axS1ubte39A+Q7kEqSPuHI/ZLZbFkd
x7w9Eo1IMaK07sYkezl1r7q0D3nTN+QvbpdKYG4BM/DfQs5cG+ws0ocAhqJHVh78
tS8a/FKNwko7nGNAqqvFK1ypiJh7swAScgG3oHKFB1IfLF9kDicCYyCazWJqG+Cd
xTjXscgzh8JjeHOy/z61uaCecNhZkW3J7qHkOeewfiH4KjXAkYfpqq52PFjyuJMC
pp8XchUR0gUEorGkLBQ4e5Uqau5WGlk0shc+fCtxoNOvdNuk/zUds51KjQq8F/yu
bMExy7apOmegpWVKgjQ5EpcM6ZVm5m2HGZVHxem2XURwAsp8t3WlCd9SlCCvchV6
DJW3R5ZSxebVkCidxoXDoqruIih6Ni/VA9gN8sFKrnBkBKxVByi510OT+O8KpVqt
ldvIneB7iXNaN0rTEjmhC9EvSsf9idI8rzCGmw/VD9aIwmRi/jIHMBweXaEhjv/7
X2sJZ9mj91yZECAV6Gkpq5N6nl6jgA/AhLdiBTBpZZ1vNnWZb40IWw4GihF5Emoz
3BRkgaUR1u0nKNtIgVBtD9a2pv5UsG4fBj1Xij3uwfHbsvOXZz0FYzpJKxEzAP0n
XglAvl9q57DUVrZfF8sLSy4f3lqom8saDFaoVeLZcExOmp+v8M09vTBDdrM/ZoPY
t/t790dnsnqW8IpxLZvX+gnOkg/Pezk7xgXI9sVcWR2pMiCZRnYIPQaT4I3gKQRu
MO/F49UGGCNRFZdIMbLt3zEBOWzavkZOjNZaElY6OjQFfOUYX95vTxcevdEyqguK
B6Pk+4U93XP44/ajGTgWjktpoP5eZDgvjp4w44vEtpvQuZh63QJBKB3j/TaflZF5
vD5kWN0EAZ5v3CahZ6b8XUNbucX/nQsgrswhdSBB8CK+WXacN4Ge8QfiYbdoE4vx
xr1bCWJrKc93OeQMnErwlusVxWiMoHr3WATYQyruitnNKbID6CuxdTDpPwFOJEDw
Wik/Y/kuzaUA9OdjFP0Hlti4QgVG+ZoM9AhQ6JsmGrmn+nAibiQFgar/yEk+yBE+
6UjBbjqrDhine6hUhoOyAZxp66qs7Mw2WdpHU3fQ2SbLvTxdrUBXCQrVXAq2+eaE
4yRG0i4YMMTfZj5uBEmcRQRosR1E+hptOzZ59ZwoXQhpusB6ZTCxxX7UcNBq/at9
y0mS9ZJOXhd9aG1bKwO//gZL0D6tZYeebfu+noyPfI2x+3itHuHoVjKuCxXggW1N
SgfXxGia6hqBJUm0ovHhJZXeafQSxq1bRc1sMP2FzvIV+gdMbrUTjM2dnHn8Yyuh
tOgbmQ+FQvDGUaFxUHAquWBs/UEp3BzmcmSFy97HjpDOl2Q5D6pOECRz4HG38LFU
E7PJvXQ/h8TgTALT3VPq2FERWy+EWUH3JspijwHw6hAp20P1fLqM1IRDKZesh2lU
3RhOv7rhuLRhwv2BFjUsjf/9Lms7ENN9GVs1YTCulBou2tAhBb1TjpONKmq99ghy
okMU38g0oRGU3MNaNnibLO+KQBO9GyABVsXxojZXJ92CdlU+TZZzQaYkT8VoFOzC
6KJ5WSXIxaESiQl1jLJIgjgRktLCV7q0DR5ANVeyV6Nk5r63M6xlLp5AU2tN+QXp
rbrR0gHU37xiLDoEMx1zFIdxK/A55wimQGpZ7SWOGrwlIduEONKQ7pzbjaSpZn9h
BBDo8SVpdE1fmaYeMGTniOaW9uwpyAoNhrMU70zdP6WBLuhsCxlQ7fw+H7W5LyY3
zkhRi9JioXDIDQyKeajDGYusuZtpvqoyV2aaijbEyA+Ha02kxotSL8dWnKXrGSfW
bfjLghxTi2s+I+RKgNdlnw+mcWExy0Hi5GKWGwrKGeH91PS/rnF2BULF1n5wdPlr
x84gQiIUmDbQAwKANwZ8OoNOSgBH8gsMRaIJoizHjmLCQGplyOtiZKEb3U7ai5+W
GZ2WMEbc15ZJhl35I69Wbn2h4MRw2ZRA3oGTxvz6lJwiW/cguV43t54KaiZ0ECvE
+M5sFRxEatSPqbfSfHhxjsDanjqHOIMZQNowR+CWoYa7XSMcZNke+4DwdUrjzkNt
Z5/8EDD+2d8vh435vEcJwLbBxVWNfqv3DgZnsrY3h3csdv177E53vkIt89ZWFior
2ZlZ6izdpAtfS5U3RdlUlZkA1Wf2bpS+hOfntSo+OBIF6MDquetIDpTw1XRcRz5f
cu8497WxzuipUhBavzsinHweCK9CBZlY0lnxPJXAHGigtAua62LYyptCi+oZLOoT
SgOs0TPzF2CXXgx0iz9geGPGlEKwasTGUrjRZG9dPAq/2wqu/66hct1EaVse1fgp
sqUnik4sLZhQUNz+4ydvYFxBFFqPF3hJNooEUEg1X4/ssHCXBhGHiWWUea9ejN/z
KwFyhc5ai36jnGbJ2gtkg1ZXwyU9t/F/fnTckkYwXEV4Q4RQwIUq78R66C/vPMig
CM8/NM70C0U4Q20Lvret9syp3CbGdXSBr7O8a98E1xoskTqndsJrkS1NeAE6PEqe
LQkLFKhUYEvHFoTURoRSeDaDLWuFF8at0g2TnTqZrxRWTBLlj8ixVmhIHnq5iC2J
URk72NmoN7gXFu1mjeOwLoSN379uAPP04H4nfxQZN612zcE6lswFyKP47KSgST7m
P+teNCeEGYAi+p/2YlOTDmCi4peFjuFYUNrFV4FVROeFKtA5LedhR949agw8pwrh
pQNYjoeiOte5wpYNTjxLFRWr3Y5lK+YDmlKjEXdTtThIqA6bzcUHxlq5YV3WlG2C
9ctaQ6JUcNkUocFNDkIXGg5/WzrUjkWZ6iUeTSjhyx94e9WYCAindlvp5n+ruXGb
qfienkuvrs3+xqqyOdknemAE+yiat6c/E2KG1goXfCsCNJChX9P01StXMBH483ID
hP7rfD1/g1axGq/Eix4ZYrQtaWuh+StcWK75ZG6R7f88fiKAtWqzqxbxELMHbVB1
yNnQ13AFRZrG9bljT+fZghAKntnfStmYqPlKfEq9cIZliLarZHkZIsUfZ893iWy4
ObCBM3yVsxJUijQGK5BagQwgRjd2xg7s6Ol46xF+9tFiTpbXl8V2hxgv6xIn67mD
+sy7p+59zA7pR3ayUdp/JC7VPSnxe1IkCcN7cD9jYG725YnK8N+kqLFP8uvJx6c/
/MJD5TQ3/AKsMa7Bkxq9DE3oXJnUUHzhxpEscIioWLlDg1ecqHlE1wXQaQEVlO6S
aDfsJTZGFL1Q/c1ZHYUJGlDry8W9ydckmknH/Atp93SHBttiZLUJpWLBFnBm6HEP
UxI6Z5ITZi6hSzAKJOfjziiPxHUNWuFy3NahMXyShKUwc0EFXouNhUxSqFFViYY+
fRiiPGEUMG88pbynULvMPai2hRcfrIkuAL0As6HlWV0vvDjHK7IQThO91l8D0E3R
EU3d7tHTWey7MXSLXWmKWBszX6pNZ8WIgfIhn1oJFyGVhrwfFrpQxrgBbXTojtAW
LegC/+aKkD0lbv/w+X5YrMmWKE/iKD26GCmIv+t6dPHF1CONqEbFVw0HdXWcU1Xm
9+ddefxHSZeP3Bp8VjwbpYOCTgZ5ZmHWNYgsP/4eYWON4usn5uzhdkvseaB7vzvl
Bn65pogAqyAwJ7naysuZlT1ZTyuEoHpONfuyzcT3oA7G5r25bzUq007BGMjQeZGQ
OMjA/A2tQVaqin2326+5N5QUaA6EQSNAHLUwUkSTlZTNYit6dK2VjOOPRTXumbGr
AOWy9ZaXVuj5jd14Hp4tXtR/+yBmAtsH3zF2CcR1FalYDFrbhELY++ePSrpC+YtY
xNJ6ABP0hZfAk4xpZ0zjW9ftQgA3gOS97/XVA5Bzbsswh19dbHLhB2TmkdWr9Hb4
RJt3i2OYwT9MtEinaGuK+l72pHTivX3ldA++w1awRxd4BQylaPyOMNmeC3u0CBzj
7W/G6bvc4vaWl4DgRLlPde+C2Q0FXjFbxHfdokdXt0dKHoqBzGvDrerQx11jNtNc
BJNMwuXHKqzNVVXb19ROFmOwkE0UiE3aHyJQ28rp9XolupwASaGYF1BDz4ZdmnyR
h7QHhY9qt9UzBiFygvBsai3cr78PpSi/DJBtHZn5YuY9CTDMaYt6qcC0hDLuFnkl
D7/7c3g8bFIW2PAd0ZSp5nQkdI9W1fVFceDmnfkPVv1eFaOIgQXWKlGdjZhUjGBH
R7uG5E+5yhKIaRDk3913yDPiDF+yCX+HYNdH6Nv1xR+CvKLMI4lQqExmMoRQiMRZ
g44ImxgasyFmv27n3sP035oS8Po8L2R8/SE9ZFeKNdQPVYURVHPDahvefmP5tPVf
eT/7PvD082xZz27k37PFj0QftP/f2ZrZIAYrsblEtULdpWXukbFXxh78HeQhZCVT
06sHv8y98aUxHdgJ+h14kheG88dpK2IzhivW1lF3TgMPkBZJrh4Yfadx3GTaNpjY
Nif3SW5oZHk5ok7my2zMnrAYJqIeks1289vizFfce8EZHxvxsUcC74LTYY0n2LUI
pAeoyb2zS/RsC+ET1tU99dpM9MEEmA91pKTVslg0NDN27J5pqTwZRlyao9IehLPz
bDA8KhAVJprf7nInqeQgD0Nd+K5/AFXnxO8ENyek4I16fzlt5iHNq5eNHdRK8+CL
LbscHSo0UB3cwbJKSkc6HMx7JJQQNsPsBi+doJa07VQvWF3Lhzcr0sDF4/DrmzRD
51mTgR0PhxWJn/rcj7PHF8NM+zjlKpNU7gemShIXfLj14RLtMDeDI1RKQAr9t3Tx
ZZDCx3JBTYc1Xi2VfHhoQaIxXYlVBEN9KLo3PdJ8mpOD4UDuLlonXKqG02dr6LD4
HET31yyVVIyQimtB5MpfNW9MaP2UvwtFnFIPd+ZzPz8nMhmrltNjU1cCq9bBfHeX
fIe9guZu+7UcrwhE8q+5P4VspS7pJvDVNy4bkgdM/AR2tSOMQ5TlqpSJ/UFiaz3G
bBm44UydF1/TmjR8B/1rR+v5MxDgUpoGRT8CnMk5HHdZnbavfF0ZESobLeqn/6aI
ME7CXjPkpSOwNU6+DsstqS3BBM2vjAyeRcjSLL/AOHnv8m1Hvj4P0YtWkGaHOMyX
rW/vko3NXdlbKpzsy/Vpew6lgZmRfnljXBMyZDuuuA6nzHTYZXDQ/nktwG934oEQ
cth77xGi/NOHzp2X0D5u4XBw+qImOHcN2uHXxfFVt7HsbUoeBZNJR2rV4lQt7QNr
v1BVIV6EUa5pnmUUfWzTr2WYBWwChLDVm6lVaAWIuDx2w23pTSEOKvg00VCUh9ih
5bx/oPdz4bxAPKU0or2iGT9u/TKM3dPUSNYzVkP79W3LwGnVe0QbFeYbz3Q48JPz
RthW6dLAs7UIItqU31pXT8Lbojio1LP3frb2mf8LIC7uHAQUtims9VhPKV1e66AT
9WpjgvCiV7tV8jZiJq5Nt1Np6ixnait40gdcG/VqzBI2nsMCRq/Mj97CPZs0lK6X
q75IjUmpcTxygs1QRlqr4QsAtZxLZreNyGqgGED1f8oEc2edquUaTVmZqFo4EYGU
4iN/ODwDBKsg8yM2OGTfMNFoeSDq/bc2Rp4ealKwYkYARxLHF+dR1HEVoDounL+e
lgIjlMT+0ytN35oyILZ+1PGVZGFBFcWC+zVsqVFLSoUuOhE2ePV/gFKPauzjWM9h
IfC0GXrC9vJ2IlsTtP3B1MkfuInGnGZe7JF0myxTLLp632lIYpFj+HifK/L3HnrO
XBhOWLEChvVCMhET5JdMIuOIQj1elmBSQ3GDtMNN4Di2IH0qXiK/xJP0tqeEwJ61
JlUt6UvfL0iYZUpMfFzzcx6LJu5ZoNCy4ZzbkRcqIDmDahK/jsXtePOa4w7nVBgV
81hOzynvMN+p75BHs/N9vOHaSM4igsaQG5U6PxiqSxkS03XDm0gMFRNzPVkAgfCf
+Lj4yuRaa+6irYmq48+jBD4UW8v5Zp2jUxjgK/QXjn1XFDVdijUtiaptSjt1gBwL
Q64Kv0s6cq/cz8nKRgPcNoNyqbY5Oyla1SJ7JgMO/tjfwvJXnKoG4p/PqdFadr84
KgS/MJbA47qpLVWs4Bl2r7JNFO16Qw83Db67p5XedV9Pg4J1hgxa9Pt/GJjX6cnB
xxlU/GY5rorowxo4V0FkzAAVdJ9tFrXGf91B59AKjgR/jRDyiJpBozlO/sS7ZLdL
5D8g+TROGA7Kfi3SoYf/V9NT0kr0SZdKX90jqxY0HHo+HIA5BvoPMR7TphT7w48z
Vk+eWOenUhvPRsSWHtCnfDYkSwr1575oWdDPIy7Tr9lHJqFngylwopHJzXUi8Mrg
RiNoCuHLuapcfT5bGS3DD3BuN3lHy8QzHZuhXGQZVVpPJX3gRWWiGzc5t/yEDBGG
+dywec4jzssfhw39LOfCVSfQQmfgxRJJo6YMCO3uh+vpU2Wgc/yYo3OQwTWPPVlI
3b//UtgldpkFo0DZoFe8/SJug98jhXPsMItUU7h0c8XR0s6AeUMzEXuUetb+dJAz
tiiUJqGIU9crXxTA+5Sy9u3iVurAh7GzG+NAEHSAB14xu7y+Hhaa5UGqShdRo6/F
+4/ZLGMBAomNUf9Tn4VwcR8Vmpgkv11b1om8RRzdY9dpCwaj/7hA9gbKQOL1JuW2
1jRMXuLYfm+UQkgX4/hSJmvTrDp1kxXhmcuI9gnSTTI9mJ8LGsutPH9x9uRLFKKN
Bc0IJdd4eGvicGShgkh7wiYh9NA4ikC9U0TX2t0onlCvzSNbNPQg0uCdMHqJYsbS
94WDLCq7P2dOCp76F9m4gQc8Eot1fMntla3YrC84O317Zbi1F1kPzMvxYxh5Sg4Q
SWx18+bjIoSdOP87YptAm/4zVGpaE40Lk9g2iC2cqHIWds35b4zzrhYjeaLYupPe
T9ul+tmBjlFGLk93SXGiM/IuWDiPVfF4rV0gw/YUFLv+wRXkKWpLoANt0C4RmzEH
alVKD4XFlTAmQyKpFI6cLTUSXj2gBJ/dfeXPJapdcmv/HtOPz8c0OauGG5KjyTk8
4gUbS0PJTUQBb9GB95UgwfWMCErha2iY6p+cYiHq2XYoyOWWHbV36p4qy7CHW0Qa
TW8l4ZBnEMSRqMrXMlgY0ZJlMdjpGR7oPmlF8TMMnnfalxEoVmYCc0DPFlqZmeM6
qFcEAI9isJWrsuCZObUeHw3jwqcF6TNvptCzRLN1jdfs4TO4ytRBnymM7OkWlUI5
WxsBUesve/T6EOGYZ48h+ZnxMv5xnd/6Yb7OTPNlMORXPiXP80GIEehri7rNVrRK
2pG/hjZO2Wt4W6KbzqX8/JUczLUEAO1zeCnzfWAMFjTD3CtxlxaZOURauZmmJfHf
QRblMeMYvZo3j0KTIkc7AH2IBNJFfqbX6CBFpNp1i6f/EyoSOlKZCbUct2zrcnBE
Qvlh/SKd3PuWgSi5UyohipmH2qUDQ/wdboBZXJExhKkODHmbmVdH3DBQZtvvaet0
iXDiXO04HKd8Lspf/mp0Kw8Bf4i5wZWgP0mGHccdd7h/IXRBqlhPN7xWQHH+5+W2
GFDcdvW6ysqo811591YgK79H9vSm9DQoo/8KC/ZMhOBKXKus4NuFBtnNjjysM62J
pxDD1jfwbGQ2xQ/Uf2U2grFGPq3f93u6kdPMMjkG+XD3xNHXJAZGc5y2ArBdgv34
/D83U6HP00lVwTk5xiBZLIYkwEffp3isDnNRMx/1qFbs2RqY1+j024MAprI/FAdv
FUOUhWOjHY4bwrTYm6g/u8xIa3l97BgPcwvtSA9PHJj2hW7l0Jn+I7f+Ywnnnwb5
WeZPGQqqVyFTX6GA+naY4Z1c1bkh1HJcePFG0ejoqGyd8vu577lfiLGAglqyI0/1
0asXDRSnTL5YqDxO0anrp224ed9qTHi6lOICqDi2HvCMRKxJQqjRA1oK+bYNwTp7
mvjbKyPbLzs80J/q+bo4nSPpmun3PxfsuM99T7tC2kUZAYFTsI5Wm3g5Z2S7IaHc
DBD1Z2+Ch+whw+aXAIeZsLIlM/a1yrHrIfzPa4vn5fr7NEJl2fajhg4NfmoY6Zv5
wLNM5tdeZqgs1sAJ3/+zP4f/W0wU0HxtK7+luVckE9Nhcmm+qiTyXQ+cX1Qkyghj
ZtL7aEoh2WUl1IgDihqQGdb16mZNgZ06Fg0mm85vo0nlc4A/Whj7+bKX319g440I
seTIfH+Q0sUbDahcVN3lcwhR/bHTrgkz/9AsEeVKBZ0IvlgKcp9vPRuMG0ih8MHY
KjNyMrujW3EZDQusm2txF64zcNHSiM7164JE6zwhVpUNo5Xm0bC/G901O/5lEnPF
EbdNrjU6gMYTSsEY9S6lgzAtHsqwP3qygGiQV42DVqQLE+9ie1+1i/mD1zfiaSqE
7jmUz8ocZQg7MmD0EEAhrrDTGZNAf5JOX616VtCeljj9lpiJx9advedKSb3a9MuL
2TKfhJau1HOvakbt/6ejLTYKgH/yXQMsK5VztkfVCIAVMFYlNNkoD5XZ05TeW0U4
r6Au5BhCgR5ym72btl6cgztk8ag5gNyNa/mdnCObtz5OOHWsLqJW8a3QUbNkEshM
A8PXOeyAZR66Gu2JwaGvC3FMXIuciHpBq8PtqjJ8PO+nIPT82RNGHEThF8rt37v+
IwT9JM+CZ1GQsXyERgoiMSk197JSHkDqal8JRp50FKE/To8tEPD/ZO7pNG9GITMH
E7XiWvSGVEqFBdaQ6WN+DWV8JmWDm2zEPTitbH5IIzO3VXCiCx1Oq1pRPWHO3+XA
XYWR9WXMXu3pqnbFfQSbL5zj0xBioMF4CSQ/ikly3tBAujqc4feM3/K4QGPijcbO
nNEu81WN8PktXe3paZ0TBEPY8Fl1tANtqDGE4EoEZo4qVAeJaYxQTzZB0+CXKSxN
j4Y57o5zopGMFajMzQY5o+w89kvXBqsRBVfYtUpE2g3LVdxDQHj9LVaF6PVgi9dG
nM52MOze/9DdivE+O8Fe9fkILj42kC3haGTI+sDPvDwTHW7TBWLPNmHgjKE+N+gb
KmHergn/zcXX9PDYRuYvDobsqi7dtUBE7Iyr+uBbdSJozavUGW5wosL5phGYQv5A
yBTy8RfWW/uO4O31ZQzSL0STbN/BazkxaSh1yAJQxGI+2tNeCJ/9/oH1sKM/qJsZ
iTPN3oAtUSzEy0ZOg3tydVo6nAbvCbhKkee71fXvwElgaeKPFWx3Ef3s0xVN3Jvh
9DBww8RYSjzlTqnx67VA3xew82IbOGuBMidpSzf1XP/5V7Fs2oYz51bPYavyxrMS
2Y10ZJXUhKpVZh7Y7PbrrjkX1eUsFWggIzOYYff+5FjKumamhMW3uMYKXBIlfcxz
xfQeYuYloIeY4CAdRtu7RYAngMj0HZNLhyHp71VtZ7aw4HrDimqe1auu91GdHGCR
o2tkJWjlVMkHaBWQaLExa2LZzHQRS0Ye7bIORWaCUSU4OAgZEKcKs7h4jtGY4eMd
s3JFndTNsXRvKZFU1E0Ry1ugOEsUJqRlLW6EP+g3o6oeULP1YqmkLcz8Ir+d1bDY
8zHM75t4oq7P/zwWzjv+fmtx/Bf8cZ1b173JOHd3d9e5P/vesEnq3ikMYTAkgecQ
XgIfZH1MneEa2T7grBMgWleQlnCH17FnPhi4oAVfwqHa5oYgULPWQkuq0vbId0uN
+Z26K1ty79fgORX7w3JIy6UKKYvufQSwDLGRv45d6/haRWI1Zst0CfdNKo6+F0rD
EdDTCCPhML2PzaxNcnemxfKNPE5/glJU63YaEY97sq6yfE68vKWT8UOKOOaAIofD
nbfxzeHAXivjf/WGPlH1xqhoVRFxp2TuBs9MkE3d+LErGvNjBV9xVsIEhFMIyZNQ
3SG88Y8yzwkW6jX0lbkZdpP0LqzN9JuibmH3Jq16eiit+O8oFkR7dGHUCvJ+0Moj
Gvds6mUAK6ar7fR7RJhOFYwlXAJfxEkxq5WkWw6JkTwTyohAOBb73V8PCNqZiJFd
x29Av+M7IfmByyUWtLIG6GyoIAxF9OL6aW1QprSxaEF6krKePshx1wtukKcgQEGz
7rIJseN+8GOvzHD9+m9GEqsQq7AsMDk3PbA51n841IWRp30AR+RaHEJuHmpCJKxz
t5r6x2xQM8PbCtnv2cN1gMEp3GAIpcxnQO4ZfJmxDVrxsrXOTpfbgYSheAbO2zVZ
7eNllayQctnKL9KXepOshXr+lTaMlfIvlbfbPCbUZIpEpFidjujP9I+e5L4CXXXl
dHKcq7cpAP5CkC8aAiZgrClafgtjMmbD0CCPhfIJr4PSt/OgTKsvmEK5I2CBH0j8
HXjcWj+ANo6EoGDxb6kw9DGckSFS1gOHY5739JAFAp9GEzNJhZHSZ1sVqYRbGFjn
QaTCkGUVvpdOuWGDb98/bMploLKjBYeezrUt5HuvxjfDZJ6Z5vCfTSSO6qbWiA5W
Y3sn1zXDhpGiu2rMHCSwEBxlclSU0WeeBl4mHTp4+MSYIg8abG6k2dDvLSq4Vlfp
eTIjx6TygR95i6bt76a4qwpoPyRZltgb9YlVZM5SOdiESSnc4SVls1+DoU2Y9sCI
QMBBFkjUAm4rAq4Q8h9CPRbVXs2y/1yGPcL+QLewQ6GNV8Vd28nGG9mNnVn4cz3v
OhGaXrXX456u1P5Z4xqVegfgQ6ma8jbDG0Hh246Rm+kOz2D+42LXO/EfMCOtmUrB
i+2accQGti14E5Nub2ujrdquruFvrJ7FfPkkA8TiTxlEL9HuJK05Ala+CbWHJfa9
kR94CajbAS8/vF8WMXX5xpJnIU1y9k7YIOEjfrn2uZq2onKXjijnX+GnezRQ6wf7
BrXUFTa5bKzN2mvhPINa8FL4iDmXGB8kzL3wKGBiwijN4fHC0RWATfhtzpS8/332
hr/A8vukHEZtf10BBB3nFf06AAsLj3rRkZHPqmo0KR7XGPdqE5NxLawjIn5tNml6
Syuu+KR6oHqrk2Fq01V3oE134i+c8P2AiiOFwRhlLZO8U5G6yAJ12W4Bp6QRQK+A
amewjgzgIZ2x2dhsrTqzcK/zRFwGekTYJn+W4hKCXCn1az9g7cK1v4+PXZx9r4yn
cu41SHBsYKrZuOyy1Nre6L50jIhszjGh8NvFUEJ+nYWXWOd/yNUFtUtD+zmNtJwN
zHpfI+vWmDVQNhr+/DwsVm6/QerJQxdxOV+P4POB3JmBdA2/0+UP9ifACXMkDSBU
MD2P1YUVN+Pj7sAdxyyYba7w36NGf6CNmUVnqmAVVhXsXF6b48gnGdKUowd0jPZv
FY4FkWFMhMiwfZ7igVd4B/4A60NuEPVHdydvnCEslGxyhpgiV5MoTq+puSa7X80x
q8uGV+u527zIbfrgY3LEr1CMuk+cAe/8C6K08ZgppPKyz30YVc6BmyQ14I2Qh8bg
7LHNO1aSDnGDnakobloHREn7mkc/PHy7XoRsKvcoD0DtnTRQJs+4rDkx9GTbB6z6
ggG5icnYRIAY8WSK6KWT2tbWZnbtcGOzdLF6OfKlKutri5o/s9v1UpyTEeJbsZoG
qNLaSUrt8HRmCxzl3hhEXfd0O4DPIPyutc4Ui0umu/v4joX2UA9uZZ7jiqecUm39
2MzepTib2exK/tYppSXNpi+bkK3hXqbVVOr+PEfDwNPJcsUUKcj6gWdyW7Tjd7qX
g/QRaeBp9Hdm+RZl8jNAeq9T0NpPUGeai0wXw8MBZu4nYcsU7xGxa1FzZTeyK2ZH
WdsOMw8Dl9q6KlxEbbKGGyrsXcQwDJZIQJ7+72KZL3mXPSeBAKVSoOEKQ0Aw1ptC
PUkf9KKHfzcZfkjaN4z8D+IUcsaB3e60XTdjvBJ6sUb+dmvoIOqJ4YbLFr5Rndq7
NlGjtUSA61atpDWR7f0GolT/K0MYwVd5cAX7/yjy0IsMg29JB+QvgmiYhrWpjjH+
K7NUT+od/WPWMMFsKQP84iXWIk4w1gfc+dcCoBcsneqAPBfzDUIUdbcj0wXoKttc
BMFBAdOWIwGP1LAGkniJgULBcfXvRY6A909csijHkF0PEEmtO4bhjoMhgCgurhRG
qGzLFSIAGIAfb1A7lZBDctUalR6cDmj0h1kuu3VF4AEWS2xmuv7yjIRx2/u2FEFa
stcZZw8MFHXrxrvh06LbjhqtlXLAZfb2N3+px+7zz9T7b2OYR11IgPfdkoYxhSJu
u40zl5SB9aQFf5u5T6jgwIsIy7spmcuS5rD1yKZDZpk4AxavbJEkcksYv18YZzPD
Eh7rjF4co4btEMPta2bOSXl5atqEyeCpDU2lLxJh5haEBEh5hioiyJQtDBB+LnIT
HfwubLwpfXF0Af/7lcsgLLZSkIE69nOD+tvcut+CuvIpUwpv4+ar0t7pZ64pXH+s
9B/9r8sOJDbl4imY31og2icsLXwfH6lXaFIbwfbGcTNOHIbohgWlYuczRoUfK1MX
4NACvnthmRU/1Ylb3DpAw/ZApdCm7iijvx6zzc25r9O0ZRPj2ocgyro9Jb4gDFWL
2qD0LAXdFnTiwefHxaQmXw1yAKCLBJomHI2ZCuNwvxm49v07M0/afR6dwnpErBZE
29jr4hZtP60f2F92VM3+hhXsjMS4bY+KXL2jxZwY/RiLDgfj/cZ715qHQf4mWjFc
Vuy1Bv/d7j9uLCPJENthaZtp7ZRXwQdRh+P3U+eHYAIKJg1DQS+bcGJjW4rjljJv
9tcWMjQfN1UF+9tZQpKETugNbjKT6CWkRe2ggJdQeTfpwJO+nx2w5kdQIwNZQfy0
1qgcRhmth2VS5qnPBSPihHUlV7ikofvj7Sfcgs6pRPsfeCT1nZEBCf5LLbzTupjB
fH+VB+fjb0BBlmMdYyNjSp+U1AnbW+gIrDExqhzlu0cYGUWHLlzNbllulaKIoZG9
55J+PpCIQvV58jDY0UJpDyqrp+z5zcaK0pv1DiGGolwYGWyYmKcP05LZGbktj4nd
EkMOmx8SeWGOXhW+RqVfb1uzZuhDEOoe/EGBGs1NyJPPBhAQiwXdT1d2uak3xAPd
1Wic91rw5Zu46rBx1MiqO7etaoy/QQ1nM5rvngDuk9jWkuLI9vgjexusZImbPRbC
EBlb0EGYHKWhSkBYte2NG1XgooVtaobbuhHH8h15gMxr1ul7n8nmwVscVochwnE2
ZJRq0wiZNB8ZSKyop6s9IP+YZcrvs35c9OXPEnSJwSZxNRFzOkdfH2zOXE0VisMd
48ZiVrqb6BufI9jTHNcLcX3IgG6/VPDCcWicCNetTotKfntqeybOgtAu3bhcHrTE
UQZfCHdc04uH4O11nKblpe8/KOuFgPs0nQnhADRrcuYMJzyYM5Ktz7SZRyQpnISd
VLSztN09D+vx3k94Y3f5pNG3ZBilEx2UhlMG1U/0jhutgUT6BMMdjpBgDhMoJQ6n
gNSxMgfka7QgyPeY6kxstWNV+V2GWc5RNpKHsAOax2jmv9w2BQYT+7vf/Oy/9ygv
8zW/DRA+pCTTTL94wA92KOWAuAXmO/6f3NWtFosVbcIh2DD+JHMUDdS7EwpT2zK3
+rl2167pH0pDq/y4OELoiLfgLEZBrUudKEOOs4O5JZMjvE401mxezzMsvZA+eR/C
wk7dcG46m5Vdo2nNmsHt4YFe+L67XaSjWjfDrM4rhhdC5jYc0tuAY+u0rFO9iKab
XVpXKeGwZFGOP6Cbk2TusD/zZny+hhR5jfhZnQT8A4A3vqN2yU4iT4m9YenfrUju
hx+ur+i4ZdrCJmJXflzfEGrjewN/ugWcevrsV99JfdTsriGRq5CFdpF4sAmsQ19a
Ub+0/hodbSqNVdgH/q3o+Rk/Qtgb4x2QKEeTLEXP6NHLA2784LPoNOaLKVsLFglS
8RwMphG1weXFOM1CvVy6XgYX8r5fP6Sf2TOQN4SbdcaNLKKki8CqItOaeBNbndi2
CUVntmok0kA2V6iNKISXZhorrmRdBNC7s3J00SaRRxmtOxWuNF5IfTiMfOYtJxI+
GxDKDR2odxPeN8B6TIlOdOjaplKH/QCVYDEPKPYeHH4CrDqElyf+wEX6cejEJVht
3rWYi4D2y8OL2vvSH3uXbmIwt0FR0wsWqjnVLU3elR6F0ZrTqitv06frMaIkO+MG
fyN9Q1/50xrAmgZ9NYH/MhU8i+gYYlSrt2zxGPNviWr/zNOc9/BGdXuXux/pdVdc
KrX9ge3X8XqQq0moNzXjmHDMWKTHBNIfjlquhKuFpezk7TqaCsBGvnUuNe2hFl7i
QznoB42esD5gPlTrjjVzV4EHb82VhGV7fE4lCH2nzm+OIMsg0UcKLpvfv3lg51lH
OdFfQqnQq9XbZVarrYe6sCJH6RsScGmzXezapEMLQnfTA6ao74168yy0N8iUk7q7
wPul51oKBv1a7dTy9EYlWtsaG6qxdGVfXENhlynf9ESaiY1u+aVT9b3t1LsQ7qxJ
6YCMV8VmXlp0GnxuTTi6C9soTPvT3J/ggxUjEthJVkc4Ih0oKpbpMLHTblp35+4J
PJtuZDaa54uvhmLZeG07I6Ve2cLusVDmuobIdWILDsO8zanZj1FlOecJ14KcstDJ
6ohRt3RpDT5VnquDlYsyOQQRZpJ2yaciInNETuvpcrAm9ouWcaBkot7A1K4GQxRU
qh9psA07ng7stkwDeH+67nxLts1D5g69ow2uvSjpueXCNpUN4ysrXzBshsvLmRA0
ylsxsiEmDDXLpjuFaO1trobxCXyfNAP5C/frFrPCOEGc9fr6ofbuBPTohWl3AiSv
3snRuarbBm7/SRXhcjiyeDqkYyx/CfMv2xosy55dhqapVV3HyTfjGrfn7ZUvoWSX
TX9sd3dT61j6LsUEL2H9RhpqQxTCTnfY3HapU7y+HvrdssNeyU8j9FozvkngJL4A
8OUSTdyfKHBHmMhXVEwVapfk/ITLRozCaUKmYabhjJH/rx7ksBeSX6M9468DiR5Y
zgNT5EaE1svT9euLfkV+uCG+Sp3QmxOv6Y5Erz+sdHFyHLvy/4Z0gurskD+rHSKG
5pgUBKFRlCn6xnVNAACOb2jER7I3BspQLEZ3L83YkVaUPcCHpl1yD/OcdyYn2kIO
Vd1Q3cqy14w5gn3qqmdAlKiJsdHaHhBILvq8CUjFpGEugzyU1eCT0zC9RnxKF3FK
hWRWkfcCFpBXaUn2z3Qw52B4uQuwLRf2M33kcF3gsikOoPBmwTjO+hZowQS+KIDI
oguhe7HlwE+18Ub6foabeRDciLXPNkqivOrkmA03JJaC9FBrivLFPaP76n0Soufx
nWA5tkx/FvYOunJwDsl5DmYEh8LiUnNGIjEKn5B9sx/qKDtCKs0xxeHjMLxn3A8J
oXH757P+SOORrxTO7T4YTk0f2QjH1gK3yYscnQ1dJQ6waEZO0L1uz/9ZH2lR916/
iYpdVFjD+4toQhgs0MXGFKC5nUWyVp5sfaeYHv7kvvPEuKuiWwL/FMTI2WDzlFJs
li5WcEahSMzgGYH5CrbB/2gxirnIvfqSgBC6nI3Nl4llYd/PWoVRpFW7jLRxXDPc
sT76/at2kWfaOksJhjsViIojNLM+Zm3j5F7ojzk3YnZBWzdbgNvlTVPaiR+wTD7Z
r+5y2KPldwx1lvMzu5PoXKsUWhywKwjTWStmP8px1JxB1yEBN9enueh+VOJdOOAg
i5FTR31coWYugci2cLxwtfXu7aiRtp2SgU6+enpJOv0HvAgUV7zpPM8fqnFnZc+5
jghPmGooT/YVkeswAQuaTG+XmvvGUHHbc4i3FStiyg6iNU4YDFyV5KdXTuDtp44E
8DfDzaLs5tJAh6+PcDfHbR8hz3/J2Y56M+DzMBCZdw2pO45/Z5fHp2+Wh56vvyZ2
AZl1Q3ax/KgKt2cvToLIFfh25xlv0foURcYZfvJH53r1fh4CWxnKwlB+RbzrYyJh
Zpq7JKKXCJRy3d4ASh7x7hNggZLed1Tu71Ly/VuLTM5MH5YS4JLtLTwGH5qc0u5d
WaBImwt8JO7rj1G48XQcA4iqgxsQx05Ig1nagjxssQ7O8Qv4l+8Zny056tLz7e4M
UjObtQ3kmJaRkPpntJ38lNphxCZyW2lbUIcWMq6fkG0O3ptNz7MZrrjABJq1keN1
kCxekMS0f+7LiCF55XnmerRrZ9HqjLgUejxtwMJjveov5w0tNBmdMguZUBNRi4nG
k4PUuX9ptlPid0pr80SmlYk3NgsgY2RA3f1ONeXniGcqyh0Tn7Sz5FDh3DT/NcNC
wKnlelaGPZ8rHtrYu42eViPNzxEcRwS9oMhSjOgHDdKwQQHtQ+aZY5w4tw5TI2bd
3POWXwcyMqnbCZBsIFT7c2SnQF/QXWpu/RpHUnruMlkBLs12QIqsa9X4s6IMcrC3
XBYcV17IaT+5edDS8vxHeaDQhwNC/AM9ioKL3g56KAjtqGWbSiXyffmGDmHetkkB
HmI+EUNIzpfh8RxqW/STKsuJyY0/Dwhodwk9UgiTyIz4NKLBWbFxW+nt0Yg9CQaJ
9JO0iCgiEJn1bEHB/q5lzSV/84Sr7Sw2DMQRbT4C/eu8R01m6rBsRQzIBd90ePTg
0c/h5oA8zYXV1AfbYsja1wlNY8LpNfZotXP5tjwA2Pi3ZvqzF0SpbpGuyYoeJKBp
yQbCgorUKZIj10iLE74sBFCk6VfZe6YVzi13bb2T0o8WbXgybEpZ1BPlQNAn8WeG
Np26ybOWAK57pSgyk4M6e7MazMcBXznE2bkBmTLKiyWeHKVuW4tIglrlIfdnuwqr
NJICoR0J4Hw4orGI6MOwh+c23Acd1F98VooIrdsdOZGT5T1/B9LKKGF6bW2brQAK
Lo+hyxclzBIlB9ssi0HaUbNVVXyzuJwAuTFF09ctL7P6rikxMIlG/PSOihUhF3oJ
N/aJOU6YEBcJb0gjdHBXimnT8HZg9na56Kaif5+8kCScLBjOMC+2P0DdfUbRLbwT
CpRoxdxHDXnOeJKnhsghbZBwQi0JOOXQzqiV39YiXJqTprJaNjkkS627UW6NC7Vc
9WtjcpZ6kLsFv4zVydubGtW0wzDYQ9qQms6xBp2910jsMVVuZjefd1oSJGJRkHcC
IIQvAAsAdlQKECp5KgfPyN3lZpD6R8uBCUlH9pDovzYrSKwCfnfLrkE8X7epVrzY
UWVPTqPFMqxrFOD9uUfIi2uY0Yvr8usYG5EcsECYdxy9crZHSxnuB+lfRw0ybJSQ
pEJgr1LHaBNgAzM9ZTCTUSuEkB3dPfIolaNldQ24SZNAytR1cFhyhIC2/HXWg8T5
Np9ZHrhd+R8VgLMAM4tUVifgZaOvIYltsBnAbni/Z28rtnRMHzUSh7RPe5mmaWtt
vFJCny/ZM0tyZbw6eoMVwurJ9BuD78SVzNwYApx8txC5P1kaM+AJnirCLqRboyOd
/UXGHjytcIpLnUC55EZEtlAa2ndxuLl1ZMbdDcz/RhfBz+jxault6bEsPaT0JNLW
BfGL3/ajarPUyb7Zk9YAVYG+z0nBIbLay3ov1L+M4H40wXWxdmDLdCxKj4yiWRJG
sCOxmLI+K+GECcG39TJ5FovJOqTiRtTSaFBZ97hx2PAjTykhfTOIhmuf+pueQtzK
crrYMWKojR77tJbEphvg6U0ykSg+I8d1eJE26Ies6Uuy2sgP4nACoE0W9gLKYIn4
KFStcNlhAoAKPyq8FEY6m5bbzu8FdMOxOZWQM5Wb5SEeBpRtgQFZKXDBxlrj/Wkw
fSRR7C+60isRSf9+8Ms9CX5rOZlIPRL6BytpjDcGBDhhbulqXCoanVxuzvgxqHjl
QzIv2CrlqvqQTtheDQACDMINUT3enmq2cmL++rpe+l1n5uE5YR/49fpjlTfZOVTq
fFpr2NKbFnWAyJmBmQZDYkhnuirv2vkNx9YydkU6w9Nr8sm5KdQS7/WTtBOOLEU3
rTG+q8DwfZ/FMuUmONHcyZeL/jL+dg0SIkIqdsuCQRgAOXRZyblzewXfw8JLHAnH
m/BAxUbq9JOYRG29Gi2Mc4pgtYp5NMv8LXCIe3oZ+Kedb8P9lINb4hMmOXPHFJGR
vajFVmQDlQVcJNr4I0ejN9j7ZK9jb6Qw52PTYcIZJ520IstfLXSNJD2lhRpWEspr
GmMlKGIXrNAbbmuYZg9UHdIw/qM4/W2CGCpfqt6+LHVOFsXsmY+gW7J8JjtnJw/t
JKSjvqvFdR7jM/fiZvoeY+fRj0O/IrrhLAvYmG3T9yYNvlaskEMgImycherw+orx
UMGJMF3XhoUuDntf9CVXblsxDwFkEJYX1a3hmz9bWDjRlXUOccNALrxs1r1Su7/O
4wH1EhSxvZD2IsXzcWszQYJEqdrx0Bvcc0chiPkfeKH1QdemANfMSB8PiG+0hcG4
U+u9usiVN/OBNAqS1X5gkioL+sIgvA3TKNezv/WBEKpdj2FDc8D5sJKT47tYW292
sxXVLOpKTwauoC1rXKrNI98xV3U2Yx72CHenVdtYZMCt3tzl6vkH2B1/JRmHMPTm
73E+xmGFPPBfnWHNY4Mkw6gRqU3Bl1sD/jt+BnQCrN0cPOvXfbJjGOJE8Dugp9XF
L1axtbz0BOwDijXvzJVW0cC3B2mkJBRzSy/4Wx561Q9OzgzpZ1ipRdg+3cXunFf3
dwgy4lByvI8mae6+fA/ezaxRsPDKwDPPzp0TM9KRFhrt3FCX9vRxqcBA6CG0sahM
suT5mrP7/YUz4M0bX9/6BxvFnSfNsNQ9HjPJOVu8WEinULU0D3TE/u9lQBO5nDSO
Xb16yvtoPN5RZqyNC5bUheTbw8B0IzTvGZ5w0EpFCuk0KmTuWyKlarFcSHaF00sb
Toqu550G8qzG8y/OtDMV+q7fDB/d/gE2AyUGjA4LS/vj0Freja2w55HbXDIuCfwH
0Kr44bq+kVFBmJAj+WrRL8h/zf/gDTAhM/gz51KnuUJ+oacEzmEXiNv1sR1cQ/ik
/+lmHMpQBBLE8h9gRp9bUdYvJY4KMIxxowVtFd/ga9YByQVRSOfeVFgX+Kk1VTLN
UTcH2NDo2u30zIwB34aPqmQmnBICP4r1pkge99MjfekgH/UeTsKCE1b2GZwR0c/K
FZe7Yb2s1sHXnbuPFGg0/dOVxJs0kOBJtNRpq4wnbiHJtkZFqa39QpPQg/HN01po
FsMPeK3LEZubkZurkG9OoDEu9p5Op0WHNhUrABMFKeWQeHwiO+cD1g+BuhfBPifP
XH2wzJABFZddT6kY5goZDd08Q7Mz9ZsI75M4liVPM7h4VbZCeD9K79wDX+bGWSEZ
s2VMmvcU1cjaAC+CLj1Vv/CMxgqNk3r47MpYU29qieveT+oTn1y4lDdS2Q5QU6jw
SZaDL4J6+KSHBUcCeGzSPFeLU66UFKZir5hybSi1V1jmjeEHIF3EewF5g1K7siBv
2TPdEUQvvfgryOgQ0z0pqRMI+CiLLiwAVg5/RaXSBcsre7EngyZopRu6ha62+hTM
uqRRjIHfToJmH9rw3q3GEscQf4dbj4fvJ1y6qLAES2BhjuQXhxV4ejDF/msEGmCD
1VIOy1GksX6ht9Lnl0Y5b6xBlV/08nboXRi0Cs7DGRpPn+sBDZpdzbS7JKn5Ras7
5bUZafyRa02FE7WPBoGtY5y/QnR6dJDaM51wM3aLpQozcWefsllinHmrn32ozbMD
LfEzswOvjsSGP4b8YmBoh2INuUmGBDL7OR3OpkUGURcRaoxvXqC0rjJ7H38D9BUJ
lI8EFdGqiYkbeE7LFYmX25Prxn6GDqux0h/55GS6tK64pbF8c8ZeevKlBXokrt0R
rmfk2Yj/0TnoF5BpYwTsWpzu7MSWUBhh9JNtk6smWxXd4FULNX/WU9/h4CgFPz7A
JuZQiDr56qMDOvdjEC65W5MGeWO7muvVIapGM+3+oquMUEyLW93VOQ26x8+a8wv+
GfIDyQAx0Q95w/UWI4RQWkBJZtH+jr1RU2tdlh1gMoc9AT3oIkbsftm3+FAdjdbA
mzLCtG4LPQVbYviZV3A6BC6ptXtcXjIqlci+06LzKfNEptOLpkg7FOfI12IQHOH3
745CnqmUOh+wE2DwodT+ScBFAp18gRyiWooHo/bD/qj6kiHdjab+1Zai/gzNrH9u
htIIqgh8zlS/GutFPKG0sPfS/PAkh4KY0SHhfog7yZPZDucaM9Ljupuzcb/vnpdM
0ln8YXpDYdAp9o+nNwqDBbALKBkeKOvvGx+MORtCRkI8aQCJ6ZWpfZlRjiNi1C1M
hoTdyo5fTDuoJkxaRuxN1ZmX9pvFAuDOMiHqSFD0QhEldznac27JCqT+MbJE5lVp
m8m0YA90eJwXvrxAxlnloSs1/64whbHdWwJmGyY/5wEBENokrLPwJj1LY+fpNruE
YeHtFjBZRInDxPL5CkeZ+4WQBvitVFs+Nf5COBS8GwlwHT2v63JNCgb63/0Vy5AA
Tod+OtvNlaXbBVcnbtdJxqhX6tvnvd3PjAn56NXaZj/zN0Jp8TGHcsDxNCexBVvG
dI+gOOZfesI9IZSEyUdDB7ZpGL5iZAp5wb33m9LHd8mTJx1NNJ5zXQh38AEgn8Xn
Nf768KeyKK4/HHVJQPjqmMEfiAAPq92+fzp5PbP1IlfNoEbSd2EK9gUAYaIpr5tS
rXTiP4Enhz0k/qPSohnF+71kzLv6g6ImgeVjsXNUT4XxV9+j8VzaiiCp/z6OWe3l
TQ0BPOe6phj7dhmHOoXNkwuiiyddjDuWPc4BUze748HMQjO3REGPg8NtulNvufjJ
LrtSQqjq1MUeQIT5VwceCZRoEru7/XFJYWFm58FMp84bN2TCW9OVX8pPdX3/pijW
6RrNeT1ERiL6otig0EETW/eve0+vRhXBDhvCGcPMM9Z8ofg8bqorBGJHzTqgnrCe
TYWCGU2nAaihVX/7yuTTdqSDQDMcXGdIjtiduJlIiBUqUw5u8M9wTHCJ0phT1ykB
8a/g9ajbYXwyS1ObTpivssEMLl1lO6BxmzqF/grwWjgNisjkr3RDrntmJ5uhRxiY
8yPpWh7s4nmHDwd2W/dh/Gds7jV8MpGrb6rU0hFYFGtrQZBBzvknz2LDbfMrivma
rrVDR4vcsxwdfxO58nRa7LD+dh/iRkL3v0bkwTeUTrLEskFV22Cx8FQ/hEJWUsB3
TWtiICJq7DiHIOuCAsEgk05ZDALYnSvSBP5smfgOQqNP5Fg/J6PPNa4TJbv6Wgpo
aRizg79cdzlouRGaEMPHbEZkEhHx9xRiKnEM0XP2BdKIOAUH0L8sXaNa58eG8Oxw
2LT4K9nVk49zNfr1rdZbbyhGqTQn8Mm3/8IoYBRiIwvuc/dTjd84kuS/SD7TOlJg
RZYDiYLsicXNcBSljclO8iU9mXCfe8XZo8tOtzfQYQwYL84Ta2o9EvbiTy9i80Fy
/McaHzzp75Z89TSmfL7greF9PU+Rp7ZGasfmbVBfkmp9WqfR4DWZyw38nkoyFNIC
qkyfeZjPqeIMJTRoNmNeSiKvzBFVcIxbqp7hUUjmOEyYY7SNz4csefrixkGHzPOX
kKBt6VjH/HccxCKyxcGCSdKCvm4MU5Zl08rRfbkZ8COO7kOUHUHsOgtRexxpqSLq
XwV18LUhZHQHbq541Giov/kjnFtXh+Q8BYFF1gS/hdurIPCgcEQGnOMQRrFllCo8
8txWVKxBu8LB5oNXnJMDWZFIEyq7+f3Kwptij7bE1S+vmqaWd0fdHYTWTFdWpAJp
IS/+B77vPnHBEfMPIoGgtofUDEyzTQ1p22Ufgc18B9kkaG/8rKsXg19vh2hMraLz
UXyQp524t2UQ/86OxTkQL+uQiuHIENNdnmU8T2YVLGuoGrOxQEzfEsWOz6Ox93+q
3KtSHqlGT8KeQKxOCvHVvnam3C5OCbuK+lAqJX1xVDdJwt97HEwtWzv7z9atxo+Q
OnW/409eJXmazYwcq2ukNTY/cNWUdC+OBXu7DpLTLI0IP8p6l9VjwPmRh8yIog8D
+qrRnlvx6GNpPD28k5v87H9sk7Zy0ZPp0MRtd2f2ZCUb5jinu8+DpHnsSufjCZBh
gRZqyzrYzQCJvXJDm14jxxoBDkLT9OcVoQcn/xoBh2ebZwQge9xUxWwJcYliNfS/
sxtglgfLz63khx+3XcWsXL3fxXxlfT0SSFwhoqvQmjYjwuKfYT9UIJVIaQHieZaZ
n2AMdsYfjJmPrKVGbal1ZZrH9q1GO7GXlZMB4oJIdUsMxbuielQO+5S5VKK6NfhE
CEm4guKIp/VW85248/OpfMj0KNXsoC5nX//dfZrrXCpAsG4yE9G1qmPT6A+ztOCd
Qk0/zE4eQ3qvmAV0s8lOoY5vrZ+3S86hwYkMHsSu/koyrgwTl5dEXoiW8j4exZUm
1Qf7NhCnDZzag84Qh1oRV79p3YaH0YjTDN1V6p/Z6NvV93nVO5BCPyU70pdAFup7
oJ9gS6jQo9aL7nG4T8gx/4FKWgRv9W4EIC1RH1bSJ0/69G/xJ64Ip+y6VfJ1CFM1
U6hw5xC43PQD4vDc8uSPsLF/+4WsJUkEvhYHQnqdXmtRRRjhFHa+xjzo8xFF9iHD
rROeylONU/3QEczd4mGVvUm7Z2dEB64zCr2NUrdCYEj7CUYRv+uKiwqOAm54Js2W
Sgvfr+aRs+UzoA3AULoNe24T/HqrA8ZDRJW+cmLIufVggoOTnPWxT9fjUl2wfOGP
kkaMGuBv3j6zoH7tGJ4le4m1LQv+3Spzzx9L96Ce/+OddlZ0UvKhY5TMPMh2FXdj
GATxVNvJXzw+bQiLBZtargiuW29BFxZVvwbAtKuDrXTRzG0qFsbVX6vRS7WyRNGr
f7e+4Ru+8Mfwd0CWn1197CQBL29cSVgx9l37INKPPJN6Eb1M8LgNAdy9Lqg2ItgW
vrXWZ9QgJnEkzAKFJ3IhORY3c3+m0PtuXb52mioL41E/xwlzNFAVjbk4J9tW8PTH
qJIAi+Ki0JnE4mEO3319S9p5tUVh49tmrjLNtB1BYD9QjpHvh3tm/ZBdUJ6NeAjY
61J/u6dmR3tq2UyzjEGxpRNOFneQVBjpBTzEiYvPhmufuVQPAXHpnXxae6A0rxfZ
f2PMULDuQNSL3EYMrgZBvpz17MvQrN9i9xE0ByJ7A6j/M8MD+EAwiFa5yfdAgNrv
7O/NONsYWT4SJj69dHveXJXrQi5gW9uks+UP9wDcybH5TK8Xt63IWv4iDkt3D+yv
XpzWeeSljbxyWoG6kko26wg0x8xdXVKRShwc3YIxdGP5fEykgMY57LxUajBiLGYj
kDaDYuwhHjdrea3gvjSkJddGn3BGxZxUab8oc3BBpGaZdlnWGwTmUDQDzRr/imqG
TeXnhm6ZDA7CysouQBcF00PZeOkfCj9ryQvdxfxsg/ECxtHBOjrVc0cjZxE4Kb0N
m24PxeO1ZhBP19ae0gh8MieNOZtOh3ij8FimaY8vpCNuDOuLJyinMCiTgg5Lmzxl
2cbJ5mNhUx3eSXq0mgtlI482QzL9KYlWokj+7ldiaE7AMtBUCKtRam5ZAH6pl8t/
8GyjYVVO/KvXudqiWumx0DfwqZRSfoK7+FZU/BiAhcHeu5jsCJD+3R1lbsw47tdV
Ju8jOUXzOp60p0MDTr3v30/OvUP6t5IhMP18Te4acu6ZP/1VHKKckA7yGXz2Hqzq
MW6jGcVQxeQv2Hy7N78wmOjSEnvXjvmKJotimF15Cqr1DKKmVHTLxQf1neSfcxI7
WvYpumarOPVTM0MNNkX/GvCDFMH7NCCrKLe7C09DBT/D/xD3rPUCHy8bG1b0Hx9Z
CNKR+s7vPDy3zmGnomCJNbSBgd8ZfTpBFFrQmbazcBVme6YQynJlRdI5Pt7szrT/
WCDCL+whguK3paLI6C38UlfCDbhsMpoOh92jPItoC2kqX4PAYXq+54rSwLbh1vkV
xHsXXZu5nHT1zwOWci7FgkR/oa0HxqmW1DNlyXqaKHJv7sB/FAnZtFL86ZwhYM6J
oJRhQtLA5xOyYo6LhoEDhMBT+uxjDwLCbAfPGaj7nUn+hYmM3IWiFVjILsid84Ti
fCIuv1/ufMYlXZlHh2kRq/sAWTmfrBylmd6eNi08c10UQsMnmMU23bAodecXICcq
FoUUeEqfxOqFDKGlShuP0gZ5XrNNCzfGkwkN7pr0mgGS0aqDcbPVcjHPiVDzcRT3
kYqMcR8LXajwxjkdlwVR93hfKWgDPpNYxPdz+UWWkiJVfL/UdDZl5LxgzSE7mwtD
Jdyih2FutWrY2Tnoug8OaBjpSbkGzhKql/GhBaZ6DDeNO5C5jT4VqlrFS13PXL3x
/B4M1C5NbfZ8YC5XYNob1Qe6ds9gkjhP8N/IV3CnYTbswr9V4rnc+JY436zV76U7
fyoW+j3zt8EtvDEntlAitk5/u2p1yvPI/SATW6h0XxtQV587peCDF22S0VoKc8Te
170WfCavLpxyLHs6BNnmFLwZqmp9bbuxJMdd6aj0oSTE15M88rF3QxfdHfga+N1U
aGJ4YSn+t3mmt9+JUAQ1SkaAFti5mitGjgqI0XgXXfsQ0fb0uDUDtoBsw/A1N8Pz
A391WLGEmnTRvet0bRzkPqtC0Jp8BVbC1xMrCArwJiZn4kxPVCmwPBQTXL9c7YFc
q5h6xB6Rk0JbYziCjUX5ydllmlfr+BujUtycDdk9VS3m3SOIGDC+i8SK/gebGX+2
Dk+S8HO6wVauqtgItY8TOIhTCVOAR2Mzci4wR1VOOp8HvB0r2YYF2uNTDBYS11vl
rzpb8D5/zL/sZRTcT0Be1Z4e+GkXAXHvz56Aw5HMvXyyIBOIq0N7U5IlZpSoWepx
8oskniAGw64Aby8DvvLADKZ/bGZMdr/Ciiir09YqZ78ax31j2DW0ZP4f4cEFEqEI
DIs1SAfvuePZezJOBVplSxaypMY+j7iHC7kYDklSg7dGmhqZtNvWBaL2bNqihyND
BF0uC8+4rAL77v3cTkv3KwGNwtDzlPY8QOZYO4pYFtT3k6NkFLzI4mn1r7GxI/8R
Ye/GHNo5bCIKN6hV2oWwiXwAQjHOU5ejS04D/Hka00RQWVkAwFv4u9yf2/KC3y4N
/7EmuT41pwMmyOH4E2ml2tmCqC5GqcTgydtp/oPB0dg7NF4ls60G6N/DzWzUPzN2
bx0NgFnuf2kjAQVkSNknbbiLOru8D6u6G75Lse3nYn+TqNguhtvsTudGgKo7Qdg9
aRuZk5/fkfnM91L7jogQb1PEojv0GuVY4i4ysaJwUbmI5atE7pS2TnSED8OK++Va
fWoutAXO/vT2LiXdWCkrHOlwMx/vZWYJYjwGM0qnWdebdl3/NsfFVxe0w/wRIrIU
C5O8wHn0EgIVPChkHJBxjokblt2DKVGgsTuH/HTb4oKTVMLltrPscQ6QNPIOKSCG
7F1mCJjGga8yiy5vqk3+ophlN8P8O3zFoUR5yW3n6vzZjVZnOZidrZfJIZBnzeHm
sVL5XlVmnMSamw52W4jVA7umXexcXA3VMAUc6VDugcLSe828pp8YNg7PNMa/4kED
JtoJQ1LaosOM2V700sxMNRIFn/frEpIJZTfhrTZ3r2z4De7vFSt+EusJrLNJuybO
WfKyAQ1Oi398V9ox4wG9lAYGibbZqAdmzfS6r5Lge38uKlJZnQUYUVAiaqUf2uAK
U7dNj0jKWCj5KJlU2LCYuzMhZRabiOUoX9F3GGgG3IGbPGY0Isr1UHt0RLl0ocF7
yReYVGllYT52194O4AFEW7XsBTNH0Gras5qmsq7pYxsI7bVDDo1JIBDNmLbU5T31
8lznDdb95Mb8j2IYwrsgU+Xf0RSeVXBY+w+QT23C2LX+2/qAzD7c9mxcZczw3uQ6
ctVVuiwLj7wEKoENz7zeY4Db136nm/l+KHUXOHEzFVcaiG61ap1nNnCeJe6p8b1J
i0n7yfbFcOYFRhSq60kynwLJK/U9DThEHND85vT1yy5Pe/5CoVpfB9k3ecZFHtZ6
/H/6fvvuXMvuzS2TN5NKKYKmt58EXyogFHMgs3IE9yL9yp9nG14JqdHGQNC2Rye1
T7Xzp8VgjWzv93Zu6Ed15E9sXkOnQlJZc1lJgedlTjLJqpNwcw8+UJ+vAOAlkBP2
GBZXdLk3M0qjMAtkN0DeguJZlGb3W1FjeFfMgcAb6CC/ROJJK+MJPg4v+OhFRblN
KYBsc1/v8eoT5HKmMN463wPshgiGTQFnVrLS9KYZK0qDSzWED/hR7VYn+hfAC013
wJ0w7+9ghpnxxHc2vX/WGUR/V7/lx/OZbmimidBMotdqhR8zrF5wB93t+wf2NU2J
pODmAFdSvsmNB9htTzk9qSwYMYEjuk4rVdjjJsfX1F11eHpawPOGEFun0AugjR/O
+9J6bWPLTuiyKCt3gsP1186cNvkzJValnBkGOhLL36v1kqtqdzRWnIkxN28WmYbO
QFFAT/x/wRv8FfKgMAKiM18PXBzIC5VMmDt7sI+otcOxvRtNiPQ40hSmbYZ/mjVy
QePz4S5MUiGIRVV2YKSoyn182YpgM2QgXUD0d74FaLpyksst+sDWbaapmVJYKWBH
DCl4PKRcRplOZ3Xv3lp78JjseU90e5bgVVTlopw9qiN5E+KzRTlLWCUW+YPBbf8F
0pMYGGx2c8sZJHKpiSbk++Miiln4UGM520B2aDiLF7JKG6nyhh52AFtKhazII/tE
klivzUhdXMCOMKktasVA6R9oGCT00WhbdA8fIeUuXYq6tVcl+JUXlmxrzxwzVxr6
cD5hY35Fe4C6TogR4lBSM+W0cZDukp5XryvRtsg6jsyPZdjY3orkIahoCDv0uZLU
bNmXU2CjDcHB8ecUpSUPF+ZZNFqahmI/duaZvAfplzKCmobCQfFqPbZDbW3qFyzQ
MXTX0IeszU0+R8b8psoAaBXB18X2zZ5KiGSUMhLXr+Jf5HHkiUp4jFTl6jhZVdvH
Yr/cdzYAFnP3W57yANGiZkJWYzO4OEh7dWLZIv90yewfAnb80ECqHfgdsRDBIepn
xruDsdGMzK3qXgAOi7FwvEaZTvBinj/brtUE2yBBSVCekcz36AdyIt/5ik/KvVq4
FclrC/5KwZJB4zFtomE6S5/5Kzin4h4Yi9pUGxB+JVLB7SREar2/hB8zT3T8P02c
VPvSwPgPRmt7O3c0iiGKG2xY0DS5uD59OfHHq8y+TYpHfePublMD1rWKQ8BUQyiU
LThQu6Qgku7xqKat0zv3mtBHBDP0hgC4wsfqutlP2BaaJgPArSvrO6N+gp9Z3siY
ILYuo5SwzjqsBM04aVIW30yRiP2eJEuV5NzfeVSlV4zRkKPpXSMYHHKbWQSKp/JE
1pZpRf3Lvvg2RrobN3R5ftrXHAY50trIzVELBmN+tZt2af6pbi7ore1fDJZSO+O8
sZ6kzWJ8CRKcysjauEraVDqCkgHMdIY/mXjFjMw0VRBYcAwUN0roAwHFNJFdgSYA
ZM8LZ9SMHNWzyHlT5wSpC1s3GadI7nhKktheGAmofwLdxdnbo9Kmr4qJIFJZBiCg
cGtOrQZmLO8inEZDZCeWye57EahIpg1I8cZwQaogmQaT+M0UgBlifQ/jgG8uUZ5P
Cx2bUOdog4c4klGl7BMMgcXdd+LG11drSaALJWHP4lkbvuR1CgBaS2Q9u8/dRoPX
j+cl35CDT23EGNwucJFXzGhyTlEjbvObP8g2TryGsH0kXwcpmxH6MKNq8pxsHUHP
20HaHImABiGUSkq8V8SRsEDsJ9NW4B4rEWY0ayHfgbsMp5JhQQwpUtUXyDQ4sEVF
+8jJdGgdun26moA3tGEdSMVJtweqA9zELMzmWfmHJO4wdX3s6BZqOW3hcxMcTKGd
2ZLAu6tOwquFNrZ8yygqWwHNTf79+6E5lU5cVvlE1vG0O5+HMHlBK9uMpINALCeK
a0dcCauTvGmaez1IteiER4zn+F5sWDTKWKMczyeq3oLwujQ3jEa04BHvAf0QXnq5
PO5OFft1UwIlYo9mtnIjVgIl4Yv1CF9i0LFiex67y3WGXYui4QwqW/hl9lVsz5IA
PyvlWsANvcLD/FRtZAsjF7Tz2OIPxsD72fEPhHAnJ0wdl95tu0QA9+KFykTbmSvn
2aKUWM4ZUqa1pTJqo5Gdfx/UBFORBKEbjeVbfe/YHpuI7UfKJNurEoYE1g5Iaava
K5SFbkoMekfCyMT4B+WgGiATCB3Z+vPrqFim0U2qW3R1q4kGQPFQNCN9CXsvHpKj
yFF0gDqLc1Mo37fLXDJoh5waCQOXzulV0xg2mI548EXmWDhgNdr21in78eGFyK6k
qTrdrXzpXr//2FQQ6tdodKtfQAZuPlpMyPd9ui/1z1M8wjSWV06xrTeKiqDZcZmQ
TYVaJMxByymyrn1rA2K0/hzm0SzKKf//h5rEEFGTZ0bMIsOibODtbV1RPKAs+RhN
Z8wttj/yHogkk0+zAZQ3Uf1ZffXJ5nn1b8EIq+6INN5queg+M/L55dBNzd+m5rYF
93q8ZU68CEEN8riLvTqz2kmdNA56v0E5Q1p59qaiooF3wHTeY4DnzMKEmL559uSB
rmrne09/l+dgrhMFfk6kE/VLVI6BxVADA9FZ3W/VCiHc4KlUKx8onRxOnbo/k3J/
BKX6xpcyq7vyardWhreodP2bpbDgtjNJO8KTpVTWFDyuLpOZMy+L9qwmEWc6ddGn
TXeax8VfZd1Ycun2xCgeYPIvo2IJaRKMOzbIwCDOusfnRETqw4iSTpAkh0oogmyB
2k1EQIq2Eqb5FWYUWwV75B5RaDay6t/QYQMD2DMVcpvuQRUDl3/O9+WIJpn6B7w8
aOFTA98ejkIAmblXZAfjcD5hseaVp4E8c0bUdSmMXIibya2ALbZFBPKT9+UYOjQy
jrj7pS2cieASaz40xwO3DnqZsvhJjgfoI5JrmGWpRpQOopkUN8XvNSijfbSTOj2r
HhXkrNdq4aMT2BSnM9VMPtw6KFSmWhuF3f/hdMIOyn+kjKpI07clxhcu714hzFmq
0lhux0xHw102S0LtWHCQcyaJOAc678IlQeIE/z11WQGxNMM8v1sgGpiaL9aPklzJ
YOQJYors1HYk0NdgXfoh6fJ0hMp0aW83wyw0uGUtoYhU8zUDEDhArhqUA5xAU+Io
8yHsvX4sqqjg21sJS0bDNMh2Gz0+ltmqyaj4UYPvR5u5ny0CKDuFQ/2mJ5Dlx7pL
aSW+unFsXneI56LtDoLg2baMgMTQsfvpw0pWATCTf2NkP4etoM/Rm0qeUkO6jWyg
ymf6T2VWKxOGrefBLyOvJ22S85hZqDE+75fro8XJv5oLeEnN66zsYKyQKoqYCM0G
no6/Fck28EOwh5WcreN1KTxtg+fgFA72+MmD4VaCvE0IvsKB+gwRQnfHGaAQYbbZ
/KTkQ5pQ0BMq9ebFnEIiSnLoHUqTmeh/Bcu6Q3VXTrBoLle7zR9DjzgCnR0XlCDh
EtGxrJl0nG1qDUl9F8yAkTHFZVxslvcR0yA4fuEe60Waxu7uw5f/jmPiZAcXu1OU
+pPCjNJ93Wgb+O958B9U5VWu6b4l0bZd0Gx2eJJZKrF4UFNqDqY2L6hZSwfoSdJz
xdK/CmlzakF03v33xmNm0tCx6iyXi3e7v4sd7mXckzp5F9AMBxcrt/zOfZuhYgjB
O8LXkE0wIdmb1+qXikgOWZ5dRb1+HYEZ1mSMmm2JSdHkq22nMZYwrY06/wmrf48a
5/myOYjvIQ3Bx0anUPy73YkjaYA6yhKE2BWtGN2f2xJrIlNJzdcBLvmccZeaj/Om
suprKa/NZu4hwwT1p4kxBKBAkAxG1DQBS8Jsy5fPHw+mzKs38zjArLyaIuYUKJHL
gn7uQfOhDQpAVcTihZewp6KMRLq2QH2i6MyDgM0MUq6iJD2z/WnEtt7zl0il4C9W
6AbjQjNOtzL1sjZIrKAJuJS9wOGm+3I3Tj745pYvPEv2Mmw3oBWe7gPpQuJyCyf3
keo115ZtI9WN0OCUmdDRxKSq6fmbmTTICc4n/77lGISEvmmHuqVj+JmrFxrehiDx
nLZpWDvg9OcoCHp4prvGIcxG5dMoFuE6Pn13DqWrJd00zCDc2Lbwnj6GXDP6imkw
1P/3FS0ke2JL13RsSDYnh7w7v23jg9IJ660fmxn7GBmPqlNVwec31EW2/11nSLa8
/0w36W/uS9cLX2XO5aXSuzHcCWfIh+r1siNhX9xTKv9eYM8B4hpUaph8Cle2QFVC
iuUTQzut6Jag+Fcj9W4m5mY5wbgTI4OSCBXXWuy03JgVH00NV+t7h6/em2CU9xDD
AP7k3gs+1BpLm6G+sXDWpcmyRaEoQZVKHdMPHbXHz0doxGNSNr+nx4fRODlu7BE1
tfhLiKYZcwgWBfLujk+aV5Eu+jNl51t+ocuWVtOH3GFPiQJYBPLi7FawE/MhkrBI
QxtWKwW7myCOtO9XiUMB0Scjtb+tulaQnEfeZQtaOTM7NZBvZ4qb8KcyS2g9aCuJ
VepZGmOQ4317PaAOXqZ7x+JAiTfmxGq1AyQOktRpwWta8qVt58vmi2JF642VNyfj
XAgBO7Nc4iNxQXJI1kJEdO87u6d2Hj0MN4KxzCt72Q26LwtShuAx8fteX9h4L4iO
yyofaRzZXpLlHeU955iIQNavhLFf+md9yEtlTXPqtSo4ncbvO8Z5zmtHcnWAKJI8
gQvQy37ktlVbTeQW+hVPHfBT24C7gqo53DrWcuz6FjdPJoUp66oG7KGDJ1PvCIzr
D2T9lkadPXvMW23dWp8wVk/jlzfc7ddJ9Yqy0hLsxKRmP2+QxonJPTZooSQpSoZw
0xFLijVMGZHYXdYxv3iSJQZfbtyR6iD82QK0k+yiN5NFG6E7KvaV71+CDLDNZj7u
LA4DHb7UF2Orcd0xyFztcoam4jqYQSOBmzeeMirgxZpOZ6oIU3kKuKhAQepUnM04
b2upyMZQlm0qauLjp2HcAMMEa74qQhTKWgxHJoEUUgSBI43bkW2peY0DWWzbvlL3
GLs6W12baeDL8nMgxY0jlc2uX1tdv47ibz//FbEe45j2zljAx5Yr/X0vu+WFiiv1
ilPuwDr5/4ENTcu4NwGfDGUvTAbs1s5BQYMKZ9mG/aZtV93/yPlQTn2Addpy9IJV
dLqDo1QZxEDYjpZvbZ3GJOoMxAB7kr/nItKnqj3VPmDhHtBeuMzSTUr1YvO0WKbd
xKU/139H+zBHtuNACoAIPotGy7or/jpJm3rovdT8pElKyv7sbwali6yAjRgdvRkq
C71k0XE7VA41bCP+GMW+0bJtt8KZJqCvO99YyhRsBZR7LDPOgr77yeEsok2jLRsl
FepJHbjl3y1I5eexFXn4kCeZwBq1XM20VV3HdJtCsKkwH6qEnnPBjW3mojqasa+Y
WQ3WPqw17UvB8lcp4tZUGtpUMay2yG1XdNLTQUakYahsaKe2dEyGN1KhlsnpzEwb
kEaR9ddX7vlOM5t+Nege+5enouybaOVLHLefMO80tg8BzkB72qkfN1jCPOjEAvGY
4a7GTLvd7dQ//XCO6Bt63fwFLCy0ggurxj+IwbbAnPjfJoGeZxKR0jJHE/8Q2xei
Jw/ys6ss6KwO+fySsDE50qOOYRMY3gF2Y/dGpIhNely9Q0kKHq9sm/EyDGAgU/gv
236LBTR9e09WSEEp4Q7gAAs5eYoeVGtELKdc3ET/QVjAzBItT4rad7+oPa/An305
Z7LmJ9oI2gh5DaOtIKOVqF4E8/H0pwdU27m38uLSR+yQ1+Se8ofkVYL6gSAv3VUB
hYAdxOGDaJCo0V+aGC2TEndSlYWUQDbT0iYyvWGqLd6giNW3F0bLPf37XVVeuB7d
rHmarLZbiHES+MbsmNh30cFZv6lFh01G46uQqAeQ5yczbcpctFIE8m0k4tP3WQ/j
d+ut+q0f5iORlfuxBLkKabQecIH41TjVMHsSVD4C8r2Jcx9rA9Gg5qbPVC+Aftq/
eda3rwv/KL1gJ/6GgWUiRtnFceyWvAae2u3ASRZfyD0f7J39Vwb11aaUHq364cvJ
GtYhadoSSbzY4ucl7nsItJ2eBYDN4Fbsolv5uY2tyawOV5OEDW432N2gnnWj8Bba
6l5Z6fnH4iq+iA/lWq+MHy7fikFlw0aK6nWos1+Ri3C2aKpp58ytdyMCCgcrkjNj
BcgoVkr7EFFRyPwr3Tgf5JFHvb+zoRNQrd0hNBvTSLPO1CboXQeRWQ0KINLjSn1p
73A90aJIuRH97Oinl7F8hJOtOExjE+GJfjssXMeUQgqZrG3bo+nThhlOB0Zqd0XH
MaBf+yuCcEM8IDNJh//HP3wOg9vtl3QDD2+dsVA5Sj3ZgI4Enbpv3X0p+s3yaPCS
Xp7YJ9D3bE0ig3UCI/Jk42+82wcEz7douBVxJhoFZNo0amg7i3/Rt58jpndcxRjM
IfrieKyhC9VVOe4L3NW+qWuhxp1h2pzAHPZAU36cAHmrGbgSWNIguvOKS1EVorTk
I4JqmCwzSDfe7025IiVkHP7ptbQywWdDEANUnvxHk+vVRMXXJxL12P4A9c9WQZ+q
HwSeVoAQC26khwbD71IQTtvsiNWcZCXzV5VGl8nhegSohK0s0jzNb/F68o0HQKey
vWwNGVnwZ2Hp2yLRpFp2Bgksxsq3nuUYfJ+ru4VcaigRrQYH9ZR5uEqvejER+JN7
xUR4K9zMxcXqqGiDgE5pzKJ+1x2XC6Up29DjL4GOaQyyvUhR6nG01vOf6CMXpjeH
N/2V/QKsvypoE5m+469QEG/4POm/hw46uoRF3oJNzqs+7zALD8iTmJ4IHj6K9H6G
JUTVvX8PpKLuvTvhd1++Bjzafvntja8kpGOQbCvkzfvkN8zvp39tko2hmgEXKNuw
V1ueiQyp+lL44jnwFbVrKqTw+lCBYA1NJ7UYU10ZP4bkWPxPqaW822ri3Lv4qgxW
PHg8RUNMMCdZ8eWtF3ojB8DpV8NawNSB40sCoRyCwpcxXPuAmG7IodBDQ8W58rZ+
0nTa9vDdkQkIHsZ3EXpSy3WDAepPfEu5FPr7oECGmtBIDeVnOh3Hg/Xz4TJYRVVC
pZFJy4EoPJY9xmfQAohtq2KijyW17zZGwyffSJeYSHuqbItcuDwS0n6YYhzds1aa
woO5iBhH3rLhTTBZCCFoAEtmEff7P96Jsg/O8TwwPIqmRXnQnwqlU+YFjQB5LikA
+pRIGY6nGtJeD/elp01IXDGLfoIjoNvGsq45f0M8XpZgKeE9oDkRd7heYogbt46V
I9hh62Yh2cxTGQUkxEL5hi69PIUa0/QSCpSDtoF0u/z9MJNq8HVFN8WmYkLesP1X
7pbKJV4I0v2ZSa4a8Qk/lm3YTmVsoo6ypyRdfwTgZCPFDfR+L9pHf2IefHph6c4u
GIXNE18CZn8be6Q8MzWvy77HQtuYRpGm+Kg8yQtgRrdz9r3oF8tsY5uL0lhOOCjN
tyPzKVoPwbxvxSg08rtfhZCxrJ2AdVHgndKpthh0y7ezeKTJnYlOux/iU6mfq/Af
PQkP1feFOWDxPAjXjPbFsQ/0lXmTaftxjIJ/6TaHnW2qo+E+vq+e7L33NkeQmPeQ
NtvaWbAiiE7Sq6iLAnTxNRAJv1Gl4oN7yLnl/Y8xg1xUN6Z8fKfU7GZ3PoGBsYjJ
YkRLohHf5GfIb4SoHGtgmYBdTb+VOgIvnHHzN5LsIEunZZeIblatU90fXn2/Fbkh
kQe68YQK3pk/xboZhglGQRLevFYfal3c/mReRD1ptzMlmUBEIXRvll4vHIEJKxFe
DsibwbAvjfLHHwy+siX5e4yBrQtcctla8N6ouPw77zbd/BF8zp1n+zdj5LGuUApH
Zj5yEW8cZEH9BXhzNQhB8t7I4kcW4L9MnytKCYC2GApaLyhO0Sl8407WJIjEyi8T
rzKfUCL5+h6/7sx1ViDo4YuijJPLfTB0Dey7O+to0u+1ZpniV13twxts2WLNLIhs
e0FZHUplIPsCQRNQQ8XCEZUI/AbjHFI88BOWpdfh/G8ApAnPGtDVZ+tRcatMWF4J
L7X7J5Z6QQp10+WlNw1MtYKmv4472xjwUxL0v9ZEyR48mFV2KnxP7lctTs6L5ZhD
HmrEdjOHtNFleIFmvQdldHxTVxOXNzS5SW80Ecu1ML49Is8dHjySx9OcfU957fI1
d7Mi/3ZbpYPVZD2ez+8sLUTP3M9wn0A9XYCSqEzAQSEc1XscVl+Jpl/udESpqEZo
r+yReSjWye3IZWcJ026ckM3UViiQU2lsV50OWNa4FynwLGox40zk0qm6LBM0H4oU
vfVO7Mvr3eFQjR3a3xEjBXKi67BucZlY+FabZooNrnopKbO4M8L+wKb5OmwnRh5J
zqoWfl3+WEys/WGHVDRsKswPbZFLUdXtUncoxzP7OPso5ywDKAspxvcreNOhx8Mi
tafMKdx3lF9DWSyGJyKdSWeCoXCZmvh/3VG8ADSVvCPPO5+Dx+ui8CJAcnOk7Qj1
m4kYf+1LCChOJySiV9EJjMT0ZkRM7H1nGRdCzt0sk1V4GaBCU1ASfkMKVV/V/hjm
ngo3RlkxKCCr5OQfhhCSQ0yI07qJYLYAu7lW5I7D69lGok0l2DA8PRSC949SHqc5
STAT+huXGlkFRWIkfmk0TkdQtEB8rp+ECEPQ3geM0xP7pp7TIX/g3IF1gqc5KT3r
e2y0eCXpEga6xECGJV6Qkg8+gUoNIY3Tn86gqd2QUBy1STVwY69U3IKLXbPNzG4v
UeLnH1lz2umBIwLEGuyXn+N5kcnjEh2HIIPAQaf/yqv/7A/LfGID4w3m3ZWFBEzA
fk8nv+P5W566RKuKb4K3DTTY/mcfeyxUgTOZBWZpTzONDxiWFJkLZtThC2KEl6EJ
pj/TtWTEKt/fm6DlA+lAQQxinv4T4QQY2RMYTP7S7i6XsvTWRNCM/CK81eU1NWup
f0/dwnoUCTLzBhmzHR9TVPrWBXB4dovwSALtT+CY59H+NUX0iTWDzRpkgXx0LQLC
ak+VsF7/1Wfz+l+FCx5TRM4FyEQUqmbYWFGZ2nsEDw3HRKltILu1DfBeAv3A0sfF
ZWUk8Spk4/K3g5TGityzqt0Hk47TQz6Xy6Fpt6UurrJbhx05ExDbsBZX22xEjlEk
0JxK+/j8sSL2rdMj1h3nmotifidcO5v/fuHtQMTdJfuvFGSgrFl/0hrF4/AfTbyt
+DqE5j2FY92ZsmmlvArNOu+ol/Ke9ke/IIWAImCIBUcPLv4i5nuSqtttkJgncapn
5ZeqwfU3jZrZiNClCnE0hy595wJU38ZU2wVeHA/Guzm8rWoymAeZoXdzUGgy+2nD
YpLervDw9psIa96siMhxhD2XLX9VdKi2UEdbzrh7+4TbhInLaC8YZbr274TUP3eL
rIkkMOmUURMotCLDE/7nWPkJkbv0ehJbl+qRqZOhn7NhslPPO2pwOtbXsW3o2wrs
lR5E339HRCBkvf5Og9HJEautMjle7eBG3fTHCDRKU18lTIlZmOBoa1OIsDrxOC38
6dKBipO0EH3OrmPOa2BroFeYzRLFktwZ2hP66WIrhhZKxv8lIil12wjOAjrI4fbp
HCSjfLr0yUxsyL1IV/IK0dvqnvxo/kREWepF2XSUhLrz4l3KN46g5ExeyGCiYa23
ov6qlvOpIZXiEu23Gk0nyeJXxcShtiPrUFOXpYegYYqI8FiAxohgz9sxfTN9di9P
swQjgS7Vf18hPjifKGozxIj1vQLPJzubKhZngEhDkj7Zr3XVCjwMdd4RgVXIwXWx
WC2+dzLSn6zEAzab8fvsmN3t+QTBdhPhuDWtcmtPL5iuixN1oCq5bG7W8HB8mObH
v3hetFSZs+F08GEoiYx9tzTRNQniR1CpjBbfsIp5lKse1Q+Tu3b+ezKJwK8UMj5q
4xYzzhppQ4NHUhV+h88JNNLYaO80YlL558WQ3zjgBnMEy47HflogzXzZfDXp3y+o
6lBEbibffyaSFvuqNvViTl1lHsnn0BRVkkbR2SOP3xMj0Bk4V3OopYCLhQ01dgW9
XaYm9p7I+Uhe82Ls8nCj6Mwa7/MEX3Y+uSrN966lyGKUgBpPl4olzvAIySy61uRO
jO52S4go+52FuDjRlIWq4D2RgiOvlqJCxknCokknW5EvE7g3b6dwHiWOnOWGS9yv
WWSdWi1vmD4ua7ApfwkA5Fu7ViARekUmxyFQmG3N1guwa3hbtANz0I+DAxb5C8IA
P+5lAg/hCNS5/eEhykU45auaCi1yFszTdKSUCU7FEmktHozmg4f7bmvOnpVvU1JK
EnzsisvCKyG4J5yqTiR4ZSYZR2f3DUUBxgZegtfde8uGPqTqzCXAdvi2uZef8w8U
pZ7SSSJdqssTjyDe2DYNyeSHVNU+tXd065PAYSuhxYgoAqp5tZKULAcyiIDhRWaZ
7tKUmqyoi3r9lRfpfwqOlTuWTUqY1NDmbllaXtetea+zJfrj46opyIPfHdCoHu5A
69IwVQajTIwpRGc1iyR77uZOOaJMeRWwvbozivm+9q4EZDbJ9Rtu36wjxlGc+sVb
K43Jvg48p3RucO1sVZ11p9iCN05DqGVLrM98PdfbDMNio5N5wMBQFec/VqTX/iEC
dXkSQwFeFhZNEb+Z4phBtcD+j5knycvnMPSotbe/UXBhvoMb7Ux0Bexu3GwLJnVC
oc7e0DsYMqP3h+JLSQsZk0FnpI9+jwEQatY3i9w5mUCRDuOcnEOqEIPqw6sUDDu5
u0LC8KUIsLS2LMEvnvc+C8H7WDrAHJc0pNGp2pKFPOKbw0CzUGXH2Q3hSkto0zrg
0MxS30rbjrWHOGrABg7UkcoXjcExBZsXM5m+o8eYqC8yIj2UCdBOlHs2x7TTyGqZ
8lYcifBAykdG+6GDqo3HMid2yf9BtPaVd27Lbng+Dk4vQIcZ0TeiFWVXaRSgDdAc
ogmJ8BnXg6Hwg8Qdna4+y22INArajru/nS1HwvQOTTmypQDigU33bodNiBCqlUNM
v8O5ZOujANvSKcW1XcJ62cUzQP9tBkQKwa8fKxElbkPDr2ULTwiV92Vc1CP4XFdh
lN8/qA2gLeaexvNNwue0uhaS/nMJLhibd4QQnUj7Xc1Y6mFa7pw16TfbSgM5+kCu
UZuEFKU79r/HJXvx1tTGxkW4hFK/s14LEVLmlOPOAceo8OoBQr1sFLZu2TDnXa7I
bOIEC8bENUcqDHPG//VN4DF0J+esqlFFlvIfw/YjF46Ycbqx6ySd6rTVjyH0SiYN
Na9UYkwHULoJ81pmBKSo599eT67vf7V2Skfer1qG1KWsOyQy6CP9qDzmZqP+otxm
pPrBL1djQWA1lZS50QzjNfDBHE8YD3n94RpsqxsJTKUkgEQnPbWCIt9GePn4GE8C
IlttZKiVhDumlqapn6MR1g6QH30whm9rwlW4GlaSfZ0CHizPmB1sg27v7MghyGPS
3AvCq4h1x7qEFltvyD4WGVt5rz2UXJLQIbu8C2SpL9I1Z6BQ5puctoAerncpr5gl
a3GNe6g0pGhpLj1jM3lxYhtR1fZj9V0gQZmqQeyMatqatwH0Cm/Vorg3boSLN5yY
CPXF/Rnfe2iQrHTtT14Cn36HEXWJQmL2WvPQ6cCVnOx01/hGatoDA29PGxvwl9Sq
uHE2wMrVyzXV3wz7XPB48hQinCYc+Mx05xeUSKOiRCcQSFWZZ5bCDzEXQkzklOBG
vQ8T8rkxAEmV3uVaIhuDIZNhj1VDDeBYoG6E+s1nU8SONy+geCoUn4WxIIhMVA5G
BfDEwDVTamuLXnQg11QPwbECh31vJCeGQ6KMP5Q/qK1hEGFg2if1Lt61nbzTwFFM
TsqeGIt2x1L1JbJ6UbhYwaMMl+S8P8RgpLndbeRBNhiXC8cVI9HmNHsrBN5K7SaA
5NY5SlGRqV5+p8uj+mBekkgKyKKyoMlcn42pwA5xAS63Y9HdXZwRKJ6xXn9PXR9N
D4F9+ECNb50bVE+bBovOTVM2wXSYRm+QaEX3s1AmJwA8bc5YPdvxdFLDVL/0yk64
sPrtnpxWeK7MP47mQ+2Hp3sCD12X21JE3Bpv8oXqG21q+QEpnnT8JM/rd3J5ea/y
Sfy2Yb7MBj3ey3XPWLZrgrvfNpPVh4cCZstLq5GQKCk/doJcQ6p/yuGyozV/dDKj
8VtK78LqgLq3/1yTHPIl1lkKVQwLJmRrMwrRHXiVGNfoayUWsGX239gEp7gsppJp
Vbg9edOq8Og3xH04h0q7vT3HZkBbyJtJKRNFCTtlY6Es5z5SJKMPwrdSRbYnUFF/
HA7yGLd9QfSFGstLm3Y4QQAIePRpb5fkYSqrLa3VnDFnza1cVxRvLrSJLGXV3u+b
fVmwRvU2wUp5jB0kRPzMEV5hUm1Z9poaIhxnKnWLX8w8nvkzt+jQhuRChzgyWksF
yUwEPL9v7pHc6ioKmt0yuwvNAa6h8eNQVnVio6ug9MQ8iH4u1Hxi1+qnZk5DK4+x
Ajl26fCuqNtVxfbAfxNZ77GP0KAIAShL5XUild0P/LBvhkbxAFhB9VcFqrPsIp5t
jv4ZEinMMG9CgqxPZ5Jb4Awj0QcFixcCRv//zNn9zw11QNnckCP5N9qEz9MSir3a
3rLGZmzinec+0m9WY08e6y33kQPXVv92kpbkbuj8KQisabpt+EKKw7zsd2wMzFaW
QEH7Tfvj+gJRPsi26uHhMRdK0QK/Qxvyv5yDYGXD0i6zURyDibEEAREfSb3IfIK0
renCnVUeR8djIolD37pNB5nZMrMD6/AHrSF0XnjeVzPmtdv+YFYe912oDtXUu8EA
3vNpbHjOGSdObgBVzHe+JVqgHJHJJCOQsMiyXp4hqYvsz4GbksCiEQFfEyO9enQ4
zVStnQL8adtCBW/yY8V5IqQpZg60e+WpEyKq5Hyjm/DGpcMH0i6u5XoSPCZTwPQW
5zHHOEaOwWG4JFML3OQBhBuWTMLisMZkyikWRRzWKTeMo6k09Kt3LQ0dIRrj73E8
S+jn92nqWr7CShB8+zYzs2HM+8pARLD8F8u74z9J1vZtTib2bIyKpuw8swNEngV1
8wD38cZgFqz3WU2EVnQvBjUsVY18VRd/sy8wG6mvA03dOYzhzrgNr5+/Pvv9hzj6
URRzke1vlUKuz7SYowkD6mEqScrnCEKrIJekJtnOrJlXCSHkiHZpA6imYBQJMNcr
4N21FOo2+TS5LsJL4kzZX0uaPZRMVyc3HZ2735S+2FSpcHXC5vheC4HCw8sPFy/e
ij//Vg6r8Sf9A0xZEpilYuCsP1B7+v5NdDxQJMzSEdI9M7V9/hLtJq96LOrM2/C5
D1Wr4xgaXMhVXZBZUjmL7QXZYJOGFBJ1PxFKfmyq/T573RamKXE0mPUStMEqJAtV
URqqqvdgmyThz9L5ZGOpSqmFmNTxAE2AF+wgs5QROlMUI4Jk44lMfgvcTgeZXaW+
tVIdmTk3cIkdqjTk6GA+bwLAiGLXWBGqm7skmIuN3byRTWh6f50uHTdsB3MCkAKL
VNcyagZbfkIMgIbIGefGheyO2dkH3y0oyEvfbGCSmIcWvXuAYMTsVCHsIRSfOQqy
xdzaYtgO042B3d/pxXrEkG4tNCum+XkkKGXRLcUejDTE6Uw6THRhlAafic+L5DgT
V5Z6kPcpmaUt8woNnNSytlQdJvxnBH/MG6syjLbKByUTf3WaxDf8UykYqNYF14Fa
saDIww14LRpKSGjiXc2l1+TYZAz5oFUgL4sxYkBvKCYVt9k26DuX9BOT6wvqXQa0
nC5DVAgBD/jpQcBH+STNBjebkaJLF5CD1uAR4x+ehyTiDiTI9lz9rkkwtCUO2tXk
xRWeSVV9Y3SsDX1lhxp7QjBvqIQehkwfyTfgfHWekBubApwf+MQg0Yt1KKzz65BA
31kCAppbbDusd1KbP9LBfI8MzVE7B2RNGE08DeL2R1VDij4Ls9wArwKvilwRFPZH
vMt/a6a0dQgoyn85ojwRuBQldCnO/8ltpmJv8l+EgZaGhK6r2kAvYpcPa4mqW1LE
b4gVoAtq5l5x3mWsu4Yn8ooBZ9vzfrfiOxv1VYdhkU9TYWsHWyRoOiUWaR8f7+N4
r0X/K3pcKZAyPWx2trCJxIsPUuiiOyJFjli/vmrd6U5ICAopaIsVysfZFrqBEswG
g70786qpNothNvvolzEl/SYKv5OilGMJhxEHYeJHnQv7FfVFHjtE3k4HZbIOw/n0
hOU//+jG6ja3kIsWrnKqCjfosq4BCa25WFiqRHw1ZH49EGQMPCxcFktd5+Px4yLq
nSOYRc186AJlXkQUWpdREGlYHnLK7S7fMwmmBVXP8o9CDa+e5T9eeWbiUs5Tgk4i
rO3it3974AlovN2TPnLc/2BiAXkjqWNSQLP3SZzuN/p8fUoRifm1jlmYjOO2bH4B
AStW/jpQUiK11Ernf9nNqkZnUmlrYHgUsru1UfqnTL8FmUyypKOOZqnAJT5JHQzP
XiWuKiL8zP8oAgF9aCGMSYd2EyZ6eTJeabLK7FjWxL+c7KZE+K9F7Q+fudN2Z2Su
UrsKieVre1PZSaGffWBOf3c/jSBS7aNSzf6kyBNHnl/KU+Tr9cb0u7NMsmyZxuZV
bfaVhF/9GnavpBRH2IzWlITfWseXewQwDIhGf/QFg2uctPFSz9vOMjpbBZ4ZpBzu
P6vr7yHEn2wy3W4nmAxpFWFJ0zCIFeufDG4/1w5IMx6o2dkn3MJ5GAcyijxGYA0S
aP3tF3B6d3ouonQqfcs8i49fw6ER8bmnTjqdrsmIChR7qNmjivmsOTXC/wtKOmHp
fPRhtpbVLKYa9VfQqtC/s4cmvfRqQ3+zKtOp7mFgwDcyLiDIcHlukey4SpoeqT3z
LEBlM2pXqNQ9c3LzlskTXRUExg57MIyV75hoklHzKebHtTOSV31psq1ewuzwt5v9
i84VKORk+un2UAPS73Fkmx8cTrcf0LqpnU8OoK/YbHQsgkkeCa8J/fIzHRlI4nNV
mfHSxJzvqN5C7vD9n4Lif+VqoT2TwmNIaMBHMM8f9+q5BBM5r2f2jsUe+DIPdvM0
iEAvZlOYPONGR7TQvGadYKfqQuYhGz48MSjGCTeDEe8P0ts+Fkpnbb6RavpQ2STf
r/5Zym0T9njS3tEkS3wObm7lUNZnjLTk2caYw7jTm8m71/0iYn78E+hXJseC7DDK
dhFTgJN3fNgXQU91FMjbuZBRelwg+E0Ujtv5ejPeunnJlox/YLW14qKJxh5uUSo7
pCrQ4MEpTE+pIB3ebK/zmd0f1niVU6FBLhex34T6vTPs6lIioiUp2aPHZHb/b1uV
0BPfdINfz+cf22QgJUquqCaot3B2JTLk8MZ2JwvaO9GogTANXQc+uuTenhYFR04X
zJjeXjm7LsLaUTl+ESMdIn5Y20MHza5RWWAv2gmA2pZvX2yyoKq2CCdY5nBwwFI8
A49mwOlBDmedm+mE7mPQ4qzujooDzINOFxN3eAIZMqvW4hEVVnAZU47/8VKSdez6
UEQrRqRPXpfYVFu7T+8iWEYX3O4MT3zGx4bOs4Vu3zl30fSeFf+iz6HGbobsUo43
stWcoo5Wcn3X89sfh6l3EG/ma0dWmy7TmZaHC6NrurPszIIihkuHeAzEuGPIxmTT
lZRp7nebeSE83pOEErU0Fl9/TGK8k7iERPPtJ33rqoW1CBQ9NT3oozdIr52GZL9y
3KhtBkivpR9vKkPo7ky+IY500r3h5RBNrma1woAGxy0wdwWCwgkaITQZk1YP02Ef
a1N9QaPO4HGvNsyYCzZww8Q+Qnb5VYd4eMeUqdLhzS9zjk+spT868/i5X7I00Jp0
BhJBbZpjDZNJphFtQbwLHVJwpUqXyYVaemHBmp+k3R0MCNNwfOMbYPiWDv/W3JM0
DvaDWbXX1TCgCsp5Qiy7GuQfSCVVLUW5TELpcsrJrI3/eyf+d/ajiR2+xyGNAbJl
zib4kkwYASvaKPsxQN0t/P0aFhc/5WA5L1abVqWcML6uA4Xn6la6PhIHU5wFKmWf
6eJCs6qdj7p45jCJAHtP2Axg8MbF5J43+3zlbuG/jzU5O2zlnZMZbe86WI0AInxn
8DqwDIQ3R//++MTgrYuht5gqQiZdqEtCKafQ7j5uHDa7o/8o4lK6Tw6c7x9WrceD
TR/NQ/Oiz3eZYWzWlotC57tNv+lLwb7wWec9XREBv3t+n4Y9mTFoOzLh3ZtmDz9i
JN/TXOep9DfTlvR55p1YuLnWCXRG1lYpxaNy45KXRitVzzZtDKNj1yHsVH0pX8lF
H2myQT9AJNtbpNrzHsljLq9uXVRo89fvJwd6tEHYUNt5fSZCSqCaYe2BzV0gMlqY
pKfD/dAUD0F1A/oE+lePLojT+a9pu1TXcD+2ojcDMxY4j7JEEaYWtXwh6lz8Av09
mJ9ZTwwYF1p5soChVw7NB6a3h64A9DaNpDbrz833dmkgNQ7+VzhvlMYFXANxa8gX
11mXFLsVIcnIjnWhnYiRoAuZ99dmIhCF+GUawDSd2xeNgQ/X4jQK+km8IitEw8pG
ObTUupBZbTSu3mN9iDDjqvEBDjA940n1tkL/F7xhnsqPNnQddPKekGU+WugNNirI
/YbeT8WiMDYJv3CN64cLhKeUlrCDnZuU2FqJxr2hJ5ypBj93y4ejJKcANuND0tmG
7glWjrudiT+7BqFHnEksAtLr4mdyyBcknEfRRtdH+/O5UjU02l7EnU4SlQL9CzY8
SKOhXYdwEoJrPHPZEfasBiyQNlQroWKansR6aXlTnBGXrLTWxfZoMSVX/EFDqx8N
+tg8UMTRHS8c8nnN3PI8ZZlsAJb8s1QQXRpyD69FW8IIX0fl1YJb1HDIJVNa+O3c
hCQzBlHxR/jVeLXjyuu6ielUHRevyXm6Rt0aC0xoqXCD+hI+l0tX4/cSkRZ+kFf4
1C6iour/HoJ9vrEYFDDYMVOhfX6D2dsEPKCpsKrJ8sksH0fmF9mkpb5D28i5CXDw
RJ7EtDRx8cv23Pz/eIuHYmcHKrIFmrv+t9TD7MNnKybsfsKRJxpL+b5re3iV3HBk
/sx1mtrj6M7tEUVb1kI52VV1dOSXCXIPU+1qLsYpbfJo9212H07fc6gusXavhEsf
ln6Yug2AbHh1j5vzsBjCnMhrZvFjhWYpQ3cddDWcHEBfTjdwTDMg52eq4pbUwtHb
oamQIddsN3jG5LQcJNmugdCcTxow+HFSBfQQ/ukCpJGxovFA4x/QFzWR4yb9I/Xs
pvDoAwV4iqNwbg6svjA1XOePoyG7OF7oO4RrQsCB1KoEuEOFo1/qQRMohKcV2zVC
0TUOyspkfoPFuInZUpVx0IPlObru4KKThA29XLH4My3lvpHxBfDBoUHGv8jh43zx
3xqyhkuv6+ClrqYaBAEpUEW9MwPUAjnECc3g6RUoESmlBioua38qXpphuJJupupA
oWQwXKxxwb0Ptp8ZBp0lgv8CJ/vuJCts0z1uMH5NS1RkjSxsD451bPRey+5pBVBe
6pr+TgXoPndboI+6AklM1RkONuBIWtt5ZYYX+9/9hMZCx+y2DvJZq1wE8MCC+rx5
MxGJ/0VmQdeOOjEaoiUPESSq6QbiszNeKIfwN3X0huAlzETTa1NYVjKTD9VSjG/O
IC5VqgCombZ5zltyIwy5Ge0wkE7CMalKYIMESyrTM0tvjCVMaBlyPEDnCUzp8ydr
T7DFUOovzaLhNwkJG3GfsYkCMo3yxI6Ty+o1PTMb+XtHmiqGjxNhIf/Q+ZqmyMW0
qcTTzlQ+837+Bv2NwYM8rOzzQgYuQVR31tl2MkDMF2To5tBMubLQxzu8Svs6V+4n
rtrCuWUsgp8nTn/ZBEK+C/W0cbA3SstCHbqTkLNq+XegavvhSigQhS0noMXkySKu
WL0auJ7MdFHudLWQIOMIHjXzUEA/D6BFfNBGVbzvc3IrE/wLdk5rINhXliIb7WXh
pcfVSIbbcceFuLDK/bDcuwhPEPw3tOv9XC4cgPOmBh40dd+O9BfPjkz8TI7slWxZ
PG0JIkV/mkTdzR2CCSqW7LvE1aDrlv9u+kcLIHohMXxpRYRZmPM3YvDaikKLzuq5
9xv3Arlace8rC44LZY6qxG/tJUWF7zHvN2d+DNIGtxmeMzpwMQRkaOdjwHFqVnK6
Nq2tWSJO4y7VHDCx03pLtcqjHAFWkikGYXroTaCbVhrc9bsD+JjCkbTL2OAAhVQe
FSklSdGVlPumULbN8yLO5RdNr1701ILWA5B/4+SgOFqaUYOx/gVub/79WTuaGOF7
rNU3PerziVlYaH+8ywZqBgnUGaFcsvIRj8hHzb6Pd4OFOAItrC18fBXNry11RCbs
x+HvNOwf0I5H1yeub7xqNwyvx6XX1HFON/PTeYcu3OTN5H0QcdyBlne8LlzB99Ad
oayFP5q28t/z5NTOcL84l+luwjpbBqsPBmVbOxa4ZKxEVDPKFgKq1/dHrLUZwVAS
fxNDlZ8FsB+0pZrh3AgoRWry+urMYYmg7bdHu2smMHDeVsKaSwW4nCzKGJ7Rq6cV
QevbLNz6+oEtDZKQVt18Ag2pglu56WBRZd2N2r5NVkWv2IK6XsY6fABDW7O0Gcfp
fs6uP7ihwp9rNy3rwMhmnIIehUmV/rFpEqvizRHX7SibOdt/HHCStCH2xY888ozO
K+mnvRSSaSefIOf6V5MUA+cwblzvRDiskwNeHQqSFV7hKyj/JARu4SXJwmk5r6/b
bBredO/T25B6b5qIi+rGWsTRLhCIAGL5Qb8fxGw+prIW/pxWaHBZokj9kFhBMS5p
qZ2je3I+NiHWKSfkF5eA08gcev1SeVqz9UejxI1EAIahcmLSklmVr8xb6JWGFnk4
oY51mZmo4Tj2IlN6tUfq3bhAAw4Y5mHT5sLtpDXK8wiLgxnfWwTDtH425qpoMQFk
QBbSmF15gl6mpEWNMQ1V8oM1f/JsqeYqhCkz+c9qEXi3LkH/+ofchG0I5BNFTOsO
t6AY/6yjHbP9z32TbuEBcokv6K9U+REsCd3K5lXTj3hmmLwWjWyb/t/hS59SE7Wv
JdsbQhS+chIWCy6w7f3HnKQJ8FIg21bnpu61TJt8NkED7PdJJ5EBfNCeTp7krxcf
H2+Tef1Akwg2zuAQW2iavgazbWC4ahUocjuAP5A3pGWUWXF5uYh6yDVSnJVVxxBm
hIBklWdIQtum1gIigNi6HB3FYrEPNuxkeJ0af4C0k+78va0aDsaOgI5tO+VKbROk
wjY7S7S/2q+H2KD/QMbjy7AIfayz7BmPmggo4FIGvcTdVef2ltIRflGzG7A62pC9
vEcyb5MamqTHldyQlLnvPb7UuavCmxxs5BnbE0FzlOjvPVwoTZoHOqh79YWR6WGa
PVdV7NqefKyGFoqVzYcWhTkZUDXSAz7ncvJi1Bzeuc2rchk9lqmOhWZnIFYKAL4F
r+an44x+R3Jo6+hPr/Mxf9+anSR90+1pVP8IYg7qaRCzrn8qFO6+wKz9cIp0lhkK
hZdFW+gS2Gh5OQuFTP/B2AGIJxY9v60LUtiFRlh5ZHZ56/jZN1+wwJhgLeG3cdq8
+Itept0HFrTz1ItjxzQ1M5jZlj2IwhM9Os7JlYs6al42xIXHR9K2PDOXr7GCJbSc
XNhkix7hXVZwo4XMvZ6z1YhJX+Rbsn8GJ0/q0H0S7laPtsRlNfHLq6xK21Nl+YS1
YtTBhMDrag8HzXHLkRCXEX1Te7wLv9nry5Mt1Tpn21sdz2/90wH0fkaY4So4L9db
U4CWmhFgPA4RIE0RkwugYn1OjfFtyzOtzkzP527GAC2jjQfO5XyWuTRCfAIUcb6x
/SWSwMKE2xhqClikkS3WR20Y7wJI9gtjJbDzoIs/BCWdrSnpJqfLGVpYEN4HDA2P
A/YSBoskPNhZGY4+ExuZd2Mkvjj/FM5NrJ7IURrnuHej1qhqdKCqofYC3P0O96FE
iGytH1ew4lTDoHO1SpQzdPRZtmlo14KEaA8cxkLduoPghjbdY7tuG7w3jiYjdzLk
4DSzeEVkOKpBbQgyO3TS51EM01ORONG27Uxk/nvM9rFNtchp3koXdB/KzuufmiND
TodO9F60fa6aLbiGf9XE3WKXJ02SRuy3PYr2ppuuiEdgsy+ViUv5CgQFd5JrP6s7
TLISqf136G/Kci46aAdZUPe7UHEwmJ+Ss/+UjZ4tVjxULP3Iu3isj+3KzCnDDrGC
gmb6shE917uaL3Hd6JELxjRKvggo9Hn5zmFK3N9gcHLQrh51FAXB1XQzX50Ewx05
rj27Ke3vCY2adwB8pj0Euz41TFj0aIvYNJ59xPSzwndtQdyHsdtuJ8/Armqrut0l
jniPQit1HOsU56Fm2T9ciCk/PFq0S7a7BklhC44zPMvilpuaE4LusFrDsuClOkyp
69ITH0qH6eMdsRb4jKEXvtsGFqCxWRPUUz2XJwJfz1q9kw7YItILypIdpbJu6jO+
EbaYx7MKE+7jZY5YM3mcPaSjZ9YsUQgdvrkZxsLmX9hMM6gD624+/tqr1JW8GmrY
/Q7DNl/pC4cULmkrdZgBBmeIRxDPYt9WA1ynETD+tELE0TUJzIATirJzRkgAhle8
G1oACo3mwMBaskwmtVozWs0Xahzfmn0tO112nczEvYcHvxKDWUz92eWqYBaKNoBK
CXtlnCytrfdeJJMw8RcxgD2lC5bOPiQovzTFoEZu9vaco2KFiPIkrspoV7K9GVuC
T3tgPEL43h9QSQZUMHBeUaMdebEOf0NcVtNISaeVQfcLZTP03/Dqy/tFMFuyRIJg
O3Ky4Fm9VpLeHrcNdkTdR0Cee4jA31731MeDsFtZLX6/a+TN0jc4/uS+on1yylOi
wo6oOgdqXs0lmw6c23WFl664euVBHgXq0SfumXcYBrOGfyLuGExu5SGjD2Eu+TQL
/FiCG771lPlrh5DqxB9pOcT879R6fPBn1iI8h6N2nWbYvxR4uFDZ4YS8blhqmnDB
/ee2xnZfguda2txHQTl3Zb51V9NzBWN7blKEaonNMeWX+mgFQHadXbxIhXACFkgO
EUwgqtJQKjGHQ45BJ3bTbToM8HAQnMOjgVgP+ly5vUBIhTszl0EoUdkTYYFZt5fw
oSjtLk9i4REst+etM7NeL8qGox3LKA6bD6gPsGgv6+fRjZwo4eueJ2WNWB4IkIhT
KzN48OXl58K+zl9FoYYp33RDRZMzb622YVtVfQNDwYjXFdRM9FNYrica6epDSmf2
Gs5jsbJnVTY01zF/iTkUxYIvz1UBofGjfwvHFqZET1PsVeFacwZwaY+D0Tdkdqy7
UUHIVYb+oCEW+zFaLnRkT7b6S0olMJkcnYIRHzUQCJz6eRTSP21WsY4vp7PmrBbz
5qo0fspaaxJZTj+uIRIs+Ff8xfgrJ5U5zUKDfNha83IKLZXuDdjqkpCghHk/J87S
RUTPQrnd+Mydb3aPak3kTein8UcFXwlpd/DdP5rrNc8kL/LfXb4tcnm0JJTt4ZAQ
3NG61OFP+7DIiUov1CMj/e0StNP49XBN5hOQPWzuBpxhegDNbgt7+Myicd1Vl15p
cYmh+JtMy+ZT31d7zveoQR6UDz2RazA9sP8aX0rMp4rjNA2/QYmnrMS3/b2XdsnQ
DDhbwwTIt0/7uO6rvtrF7duzQCzlsKoMk9l4GChw9ggcH/RT42LpavJbMWOy5LF+
FXErydleOf7385NlzHpKebzI9MBL5Y6lKGuWB1226RMwNIwkHuw8MahDoUW2KhtA
H3WBvxrM5V12/aNok0UdOCj0EqUJfJwhCpDkcvSCss1SDgKJM8kgMcyw6LLOE6lr
8F1YJO7aLIc8HJlFdL9CmJ9Qpof4PmzwnhrFCksAA2Nw1+AePVWG5M6KO2oUeuGr
ygZ59Ywg0E/imCOTbDhlmX6dFoBLiy9CNLC/XLyvnEPu5i48DVyRcfyrVE8z2zJ1
B2damp0ElUB2p3em5HoGjMY46SVassXpUuTy7nCTafVfp62Sarq63GWPR6CtaFX3
NxEmlofhTL8IHDs5w55vr0TN/bfH9yhfGNVsoHJVFR4+7lhFv23MfXO7v4ar54yH
+csSUH9xv/EEH9y2IP2wM1/bg95a6rs7NitZTRo6MJ0U+iU60Xw29Vj7Q8czxARL
jtmfviN0tZZIvEgWeB8dsYA7e9gp3cnMo/3mHTXJFM7W96oVNdDeGaDNjGi2kVi/
cbC9jYJGFNEXQtRNJhTw4GJIRpA265oqeUkTaxL/cKAGl+XAU0E587pEtCtWoCPr
akJV0xIhW1Mbv9A/by4+ldadYdh1yiQMRQ64Fz3J+661hDiFo8bXKC/RDXSkPJXz
xx9lSdgTXXeoC86UT9qaeOm669CzVzmQKsseD76MKx07uXuiKgQlvp8N3sWJPyQS
+mk/iCDT5MaGfLZ+FelHijnarB2bFSkfQ9D2oA6X6jxT87Tzm+8gnmgO10EujXKo
ilp1qpotzQwt5hDMKb2gkdL192kg2HhW9zjTp1s57xmS+3eQfw6yZyPP0RQGUGY5
YMB4E5LliHpk0LlLesnQzXruzV3s7FjDiarVkFc0q/y7g1pc6CvRJlY6OvqQ740p
2jzhJBLouUiaKIyfib55TGcsNge9mzPZn3O/N4dgWpShvwXGZofm7aD2pIc8qef2
uvsfP2gDaragJcPzDojgjRykbzT/Gzpl5/4D9VjXsJFF7FBC+KNNtGGAnSt3egC4
3U2RDrFXvbBqOlLhSbUGvlDRR8+W/o5UlL9rvT9d92dAWD7p+QHklEIwU9YBCWl3
0+WPFklLx9CboqPve1wPOee3HW2EmJjuCjNjwP1PF4DfVGEr29YIr7pXCY7MwNpV
Eq46MlMCsC795lgMOpzxXYNHRRI0hOtx3B7OSYyzVraSNHJ1kOpH9duAvUSFb2ND
BHBUDD1ou7tfOAx1394UJuox1y5GBV57a+Q/sCN4jNZ60LhOHQZtlps5TcC66cy/
2cpvqD0L8JWZ6b/r0Zqxc4gvnixYPvEOCew0BnQhnCK36gFOX5RvosCye/wGpDsf
srALk/rRy15BMJC69fZCgRtHihv0eiRSU+NXiNGa3Ab8KAFa2axL2driiGVb4saq
ng7q3iXLubuvQnHsQR8K9YggyLTFkvf8gKSz7qB6EQccOmSnzt/BIJNgzInTaicN
fCoJPUjnYLkEpHa/p+h0hJmvZWBwaEisQXt/D+m/4ZgM6tZNRzj6J83p8BbM0Q/V
Sc4WBhtoqIcmU8NM6Smn4rmMe2QF8WuGv8YXbOT6tWB5TGK/LJPUAAkMMZU8Iz7g
iDDorz251lbwRGylEaXucsm49kfYj2dhOJcOeYB5RWEkiHWFFXtvLI9/XNDQtzKC
wFx0YJNsqHva77fNVloe33dhCOverYIe+FHpViBEiOtdCBpAvucFsSve4f85cbEr
ooacFWDRrwxV/81vdHn/vhfWOKCg9AZDCOOE9UGEMxg1lGE+h8mTAHCN9MPnF9Rg
bgWc6KIht+ezALZ0fc/ncEGcIFNAjsaWeO+O9reKjuV7B4xN3Qyb4EP+LdsDyok2
hy1chUw/NtGqqZBPb7+nmDeUHtchFN0yetZTQ/GGqHZlDRInB6m+oWaLqRi/9z0K
Z+qwMzUaLsZNo05CmC0w2lo2X02fAv0nEUtEGsJZFhs/OrdRrbewmemZb/79z4k6
DjA73r6mhzhjSgI257sngGlhvmK/a9/61NoB1bvBa5/hA/HHvVqelugggMuGWFZ/
mNYG1Qvh2ylTmvV7C1nWtJoCRrn4A7tJWpLQP+ZOc/p1Qp0NX8bFD/pR8HYiSjqw
LrvH9k92b63NwbAgd/Tu8UJGMPH0yiasz7G+h89LMIrKSQa2V+4Ryghugh3mGRqQ
P5eTiSIaoZCM2aiiz6U4IVRRo8DV7x9xzZaUwrhqieQDxMruInmIbBB/HcwHfWnU
5Ru00vd5l4zjaM2xmQs63+u+Dksvutlo379lR2Dj0AIXyQdCrWvyU8ruBCTT+Sf1
jatpOiCFnAAIsnaQGoHRLcOAr7pzr/2NLI5m7W/psJ2P1UhNKvNGAxqSWrHrnAd7
36qGPAEyx1buLUgeAWV9HWSZaPDUw3nd/YnP5fg690oGX6ZwqglwXmf6Ca8M2rhD
5g3C7bmCK7Vzx4Os4nJcgorHimtC3vMFSWQP9ULEDU12rjwPTpgx+vuTaIDpGubI
tz84GZRW0qY9eSrD+KgVQAd/mTsPT/O68WUHwISSaEy5d6Tlj/wJZ09dgkrgtN8g
MvvdNHMr8sGR0ocNPjKTGDuGE4pVk9C+BkjYG//Qm1cChw/JknYUrQw0ZH96JBie
NDH3ncXJq5K4683G1lrNV5JElsQxPZojhrfoC+sePo8Kn5Xw9h+4DK/4yU0yRNJf
T2zGU21Ti2BgQ9Ckyc5WMZrppk+5hupMQgm1U3PDS74oNzO44x/S5JmX5S/38HAA
fOmar5dqp0i5Yy33/713woCNTuD8NUXNDs4PzYjmwAI4RMEN2ygsyvFhLp3eFQn4
eOLPM2bMVMomA73REFf+ouBjRp/Bz5lFHxnNPYpJRYIxKGdLacKQ/bkz6pah9GUS
bUImttqjIahbrqnRua7UhpJV4mdl6Td9mMLQu79etvv2/A7dYdXDCFHbR1/7DSEm
s6/RGQKiBA1XCQ+oxwDtpdor+jaJzA05LOvu7Aua3A7KyY5Iwacr9p3A3MmeLa5E
WqIktyaJtl7PHWXlZlReC1Hrs/MUUWU3IE1Bl65/Zbzh0vZZH3aJIOVz4kiVI5JT
ocaziu+1S4RCjZGJDNTFmTgXndZFl5pQuL18PkLCIV31E2awnDX8C2k0vE/hFbYY
hJzUHkfltb/b/3AESU/2aXKRu0nxTClccnJpTMNaxoRcmKeEBF4sFqw4QOBLDRaw
1QiKXMQGNK05A4Z00WjEjP4DHdSSvN5zx5u/mHIBu85D/H5tK8gguo9qp58FMb5v
m71FAvOtnbqITK7E2aW8wq9fZEqWQ2UTn9/C2THPrV/hbGguWtiSFAnG2eEBu1oc
/z4oNRwaLQf3kPDhpNPyu0qvM+u7YrF6Zbaw2Pz1GoR0qEtIlyqiarnEIhB5ulCQ
j8ZzEt8XIbDNc5+7Bl3s670rcjunRA/lEDsJtFVx2JjyX4htgQ7N5g8miCvsn7/U
qrqxStfX7VXXGvCroFHTXHHm4dJTYZYBphfAqRSvKUpEDARfN7WW1IN5Q6/Fmv2r
BCxX0UQv3I0/Xv4wBoFLjrAd0lzrYmCAm5cIIuS/0gdQzZ0SUQ2Q/TiI6BnH0KC8
7hnPJeuowe7OMyhjgGbMTfOOQPoDJ3lnzpJQHGU2b0dMPVmMRD6wxDVMqNpu4bLd
p7+FDpVJSqDW1yusQbn6LHQ6jKXej8qKYrh/6YSBJkpqG/V9J7hHfHC4S4oKwnwN
+atZKT1ZtK3jJ0JboYpolyTWTxjQfdeA6tutr1bWK+aEjr3PaL3PaXlhmNCKETTP
ywY9ew9Ngvy2DJVu4x/3zkREx91fzcn9ScfLJ9vF4BeiRPPRkDnRHWKweFrhHuqr
pCHoHhA1ZdOeEaqnFWpxaKwnhgzDsbuzckJtPIWtaLDKLKV+A8ryDxvSe1jh3+Z+
uaroDojN9KlSTFq5w6i7Mx1Qjosl5ymw6oWtWdSOM2fAQay4aG8TimX1SB/Uyz1u
N9fjEjdUlLTYOr6G+lGO1HoQSuS3g/UwtcXFJw4QKvfuFma7U15SwwllDTTSmerK
V09MCqhcLCU3ZvlYJhQfA0oXXmOCCCd3/o0zGqCSrMMlEcJxr+D5W5PatP/Bg+P3
E8sEMqHfGK/rRb9oEj8hyVuZuWXzdZydbnv1op4FNcsSgxbdH0vqhNZLLvO2zrgl
3L5XXRAXmxKPaUTqWX/1ZC2KDZwnvvvahDISmyI7eRehSVODkIAHJlO/6YcWbQRP
uc/v62ti+3Z2u1XjBTH1Q1qck1E+amDPRBPDwa1Jbg49y0nabSKvGMEm/tb9SMIU
3V97I22zf7KsrF/0vtjpvGtlZPvtpsoLledn0Vj+HMJp2NAPE2RuCAPt+hpM9tpb
7RLmAL1zxThzVL5yHEojC85lhaIqPKdafNKwgBOUZO6up45XUagESsyr5T7F9X26
WRIR1aLBvOTW2H95ZxaVcLh09ZKUi4078j/UaNHyesi87s4bQBO/5+ieLMv+hFzI
dZ84Ypnt1zj5Ce9iv+Fxxe3H5uAzbspNwRNJzTPPQdDH8xhxt3Ey8Wdh+us92VCA
IrJtKhvIcIWqgeqpTN4A2iKP0dCpUFTMViA8RIStNAUcSBrXfFhsk1evOE2+Lvzp
GUDzAVw3iAGVDACKjvzVtdrN1qDwnK+oGAY15kBWYjv8EIJFhnRsQAhAcRybDH6d
mtFFot3QaPcoQInUAr0dIyTlYlBO4xQDv51/hLP1uO8KQzv3rcGU6P758qAYiuDu
iDuBUvDa+wekt6jYE90/Lbdn7fscwOqTOa+RJW5omctfCIWuDLhzCPvgZ5n9LtUe
U+3h9ajKQYBYRS70tWTSF46qC/auKFdr9kbdP1wbeys8VTRk2HNQ50ZayA3vzdU7
cqdOfXMWefHiN9h1vlrVPwTfFudpm4ifC1OWtwpltfjKLl/irJlivwG8PZJ5YK/F
ffHHzV1DVsxrlJT5rZgsBAHmyQcZuxE4Wec3JRhG8u9KWElDtcZBemHazNanfix5
x58GfVz7jWOls+fbgCSv2n7Yy2Sq1wjI9xLJL3tNYVhNVugq0b4wbhK5P/SMtuLK
5lIYQhDAeo/QDJV1egu0kDljaEbWaVGHCi/oGZMubiS7mb/cdE86kC8r72TU3IHg
/iz5dJZ/fbZ6pu8jPszF6sErKrX8Nh08KqOqH1Tmb5K74lUpGJoRHlt71juxDWvS
0EgeG+SEiMZcL5wkcXnhZiRoBmB8mx7xCJ8O54FaHBDRQxp7zYVbEC7vg5S9jBSY
Bya0YENehT04VcQIshH7245WIVxGdhXeJmncKtYlfJaH0NFVHPEOldb0I9OuyCCt
lMfBZDNr/0uV85+RwOVhi7tXgPZd8HvJ2SEk+adC/CTjDawm4zurdJZ6NwIU+kOt
5UuBszhJK82pykkh/Dcx/8dbWgW1KRnxPjRiw8VZjptfwJq9wlORTE4dP/KfnyeK
uKIXRGPG0+ITCznkjQ262eNZNBS/kUSHSJsLBeuVHmBGsWg7LvR/W9IJYpeb9Nm4
blzBS0pkS49H7xBDtl6/CnNbGpoI5FRRovg7cUI30rlrgQMh8uaj1qJ3g8llBGX+
AeXKnCCAEOGKcOsE5XtVjeWoHZxCOkSIZDJuF08OU1Bbowp62kH43JuGZK+ban6u
jDf4ktN5hA3DrbMczlpyTHgkKjM6lUr0BkzTRLl1amHOHa4nr/v5raa4xgOcVWYd
3hUxf1zhlnDvXgYuG3Z3fo1Q2Ts1PQ6EUf9y9tI4OAaM+WvC0mt+L9uGM2INhRRm
wNTTc6tHUd9MCUHvPrJtyTULcRAbRiyf9H2lU8H+xaRrCwDYFcOiEsm8rDnWZUeI
+uZElQ1nwS1g0Jnj8H6yeMJREbRYTi3nqxVntj9oYvDd5JvZM8pReMzn19FKY/1l
e0ccHXJ81dICYCpkkcVfjboFhlbBKhJTGaso9IK0oJU0FVkdGhkiM6DhfpEJsBd4
JjFlOcjCgLMNeFXgAumnl7R7pg7b4qV0nskbMoYrSJpn98rstm17bWWKr2eICZQa
54DMLwWwqnh0njeaMVKOEdoVJGQw1k6TWHYNq4iUUgfFIU9Cxs7LVFpGblYskwqK
fxsbVvWJzMn0YU+Lm54n5GcTtYWiNUUzz2eMe1xYtX4KoFql778TaQ+9frLkEWg/
8zb0D9+vqGChK9fLRDXj6zwuaFOBJ6walYME6+300FoySCxcM5QaDFa1kffK7ByP
CZV71H4p/XmogaHFy4PjFeG9LYdAEbK9LIy5qkG48ncoXV2b4Kh5cGGqdI03IzmY
bpEB07wFvN2mrda4dMAdlDYIxDpCyAMIquUv8eEvqNQwBLHrbGPUgdVveB7+i0UX
/tg3w0Y0hm3i2MBXGRFs+R0hamtL+P3mLmR4+GxMWpbr/orVLn/gXYq477Pyv4mR
t4Ql97vlHpJ6ZCMjLPGxlUJG2Opkw9jKDq5eTbzZ64UUVtxjvwYA8nNNJQQVKUzG
SuRR5hpyOt4q2+overmIzB0kpPZpwdL92DZU1r8KT3+HF9v8EfYDB4/U5Pkep5j5
Go9Oc5NojLGh95RNs6bv8Y4brKLDAUENDGYjTjJV9beA85pyYSbYO8nXWmM6oMxs
DZiTlVBOK4AKUulP99z3W8h9+MmU4UOTrchkeM2AgNzCT1QC1K6q0Darpa/Qpcz5
niEuhmDU77MHZ4pUBMb1Y6lddHNMfvsEPfhAX31FxcBUVLzcbq3DDqO0rVNorAdZ
LzeeUrlN7gV0cCw5ccgWb6GRaX9WUukVB0w+vbpEKX461EaHVSO4UBIRFySjUuzq
1Bhv/J9Pt/qnIOsrNnnZggIxEWoYuJ+pfV3miINpmeDnTSGslZVOd7X+QQegQqb4
0tSuViv/PZ8cKVgM/cS49X1i37BiDf36IX7fhS4xXcWp6pQqO9AVEY7sdXtogi9q
YVycFBPbmXwyRjK+mGMdnKdHjWUpeFe9PuL9zLR5oK7rQnWVONx7xfzkDDi/ntc9
3xtfXqntjuVH98fmocAc3Iy8/qjfKh6/3RQjnXyWbmWa8cZF3jguOCGM4uQBRppZ
Yb5mKPbKCoWrfaVxk2YDSaVvcUj1dkjaqwrA4ZicaZjE+ejMCdNs7DfQ5oqGCpgn
Gi9XeNp/8J2yAveSJADLgWMhgp+SB2ru0vWm/mOeqkE+FPp39mEiGb+B+dO6ImSR
LPmvmd1Gt/MdRvjBFYhDk6IHO7A4GUqksqP1VWyrJxGfTAPY5tqNnT0MbKvPqYJ5
wuEYKaMdTsWvGa/UNyGPm6galot4dz1Ak7AHH4Oh+ttGHik5kHGbc0A/5mTB7UiO
O9wIYnwjWffMFTIRZ7ulaWjVS8VvmkOfHNr1L29dveBpRqjlF97Z1RnG6XAjeceP
c5zwrQUgtL/V8lE7vqw3lfsFsAJUnmFcqseHl/hZN1S40uPS2X03CtSUFgcNg8yy
EIanqRQ1ieazC/hEmYuc13sHb25S0bMVeNQbUhaMlWrtwrDpw+w4PiJChpWlQ8BV
VzBboexALl5cJsL5ISbJSZAzuCerFpTI+4ZmwVPWD7kvz9FRpHF8G8sS/VQJyMcc
Yc6U4D2btIO3SGphP8a4fJ4SEPmz/uFYUbmC2WGsQ0X6Pt/u2J6NAZMKuZ1b6c4U
uImBRkQWAGUZI70FbAu5vufrFXpoupL5duqRmT3Rb3OS+x6lCYF0v7Mk8RxyDpCI
ugheG5fOfUY3w/+vEIuef48CJdQTvOHnmie/EQwsDkY7VPwUdfPXMX7qoCBpli4p
/Is3asA4EDSxPkuYYFew/tXSLR4rH4aENTVycaQR5+kKmaCe3OYYqZbYUi4xSsvq
dy6evFsN9dX1SFKzNHdFvcdIa3USqTG2eQYZeyo+B+Cm5v1ICb6hyhsnIUHgkM2o
AGO3WH02lZu8gIdKQE32n6fQQMtRywbsIbe7awZ1afSB+Adwhktg4w06hYA3NVNP
TNqPx12mOwx6HoiW/MauyutMtZza9diXxzN5bqdv0XsWDF23mDLC48ygt8KpuZrK
P/KNYCpnPj0T0NUc+8STGqhYGZ4sw8QUEhhAf7ZbFsR+q4Z302WAty5YCSWOMJv9
/h6G3M7V0ZeRdwSeEWbJKjjJtT9Ek78WVUUxNvZtrQYZnXlnW48Y2u+GxE+SWp+x
w4PtvnxkeZnmQuf0FSzp20yb1MQofNwGz3yj36wjCIyiA4BmhvLg8Bq/WZZbhyZt
To/GlH1FKoQ63aFsh2Gef6N1JqU6apkDyJfVZ29fgLvdZwgrtJw3nOLygGAlUDV0
BrnbBTr1ACjMu3HmWjoInNivX+uvEB/oa3eYYqwnfFTpFJFl6r3/pFk1EoEprps/
8sPjQ7eIcggU24BYmoGsuoHdx7VE3Ff9t6dysfOSHm4BDHqrVeMNqn65SQMTJJuz
5/p15KYxYP5FeF3TH0rVTtfELdNC0b80Mk2Ud2+0mbzfyczsFkqz42cBWgxD0mrJ
uJIdlj2v7m3DkWrFEQnUjnlHK3euFAdmR2+BZ5EPqpfvP4ILLnTWwqgWYd479vLa
iSNBSyS4ZC3vtpRPekznUfE6XV3Tpda+7jOPNin9dKNoWtR6hy89qFNDA5nG2VxM
NGBPYdPBv1YkgAB5ap3H+G54gdj/AbdcNYqGZEfXTErLHYJjEJiqiIXL/bC0KYJV
1G0DsbS10I53SNPfElBa+cKblir7IM+Hkh2W23apON/yZHZJ8PWDuI7S57dETN5g
6mTCAg0q2BFT8S7RcqwsEf+Zd4zT520GycRJb9sDDbwNPd4bEUkd0cIn2hocFRY1
IrEn1L88ZRBYiIE43WXKrVz9FT5mYEZbTonuPlLWwakhlPvfTRZIARinMiotUk3p
8QBokgzKb98XHKlQPBnIf7iqIZjIJtkPoIECIlspVPDbof5oh3AZlEgRNjC1cC7l
e/4KaZa7nOhTcuiHFeBqtHd0/kPcXkMoUCmNExxLzco3lXd+j2B+PJlI3QW9KYJG
0KCI/4VlkRUg4keGlMib4rVxAGzpq+xP5VcwtbFPegxgqsq8696E1DgzUMwatlSo
K7FzjidhgOnBQPcXmOJ8xmrsqNGN8Q6TZDdOib2bkT+sMpagKXQznyc113opawUP
tf+C4b2cydfLuGSqH23kkq8jZhFRg8b5C1osz7VxGZE1ZdQhqxA4atuks+gJttMR
aG8nxwg1/6pCeZrEK5VfyrfGL0xhzg6OH7vRpxqNgaF2BRaO7WWG48JvOzYH+fw7
DErUi0rvBL4MaEAyBZAKmv2Oqof8X0jAYG58EF8JIdbnMq6gJ3RHwJYzJzl5ceU7
nGcJiMFVfCPpCLq+623zPAYdibNlpTCzavB6etvLZJI9pdZao7Za3E93upzkOTwM
zBZu4T/wEHP5hW54heTMOYm1OWBfeRQfzGDVOxefbLOOx0ciySA+P/vuO0oNj8PD
5xyn1BDtC+WWd2eSprBwpvUYwZCpzR92w44Y/ff63wARXZKMjZelnVGLzEsDVYtr
HDXu+Uz5MevIw4LiLTLfApC0VZeFmj7S3Fip8PUbbLVkIfdIwtNH+7n9ISRnuREv
dZlIN9SwHZSFFMp3jbVUD5M8TV1/z3bH4acvSj9qiF7wsePLeZJ04nPeB8qfFUW1
mr5xqeXM3zFsxsBDOgswRIaLNem7MrkSh+W2cBFokDv0csrIiW9Ck/JN+xhYbdvI
j5mQLIy1z6vL/ExjjuOHfETTnTUNW7zmk/nO8ZCUOhg+wEvrb6UVW13Guyf07FCk
VnbDKkLBFUoQPSIgKUm2EwxSlpsbCaifhpuGXItXBH0CSx2AeB6+Q+OUeEZsgYUB
8lZxhp+OOYE1R3Nq2u8Z/fQN16ItzaLIZPa4nxyy6i0EltB1Y1vtMGc0nvitbuu9
NMKOXr6M9qyRvI+82HkE2EX2RqU1/j7UDhPOOcrHD7mLRUGJvXrGN63tYk+2WQQE
ABa8KOJHesT7tgaAoTPSRs0RKKLNlr6U2FQUh+ReTwuWRDCgl8l50y+dzdVxefd+
3Rwe+vs4Ghzri+5ymaK72dA74dlF+1+DxCnuJpwjrAp8YoFkIzqCJ8FMA4uv6jxU
O5hFSgiLgUbs1WBX1+sDwvGcO5QIRHw2UV8m0fZTAbX8jlSDKJM5/ckwobuySAHk
rYIMWqgd+AyGRSE/yXckCVAeTfN0mjvpW9mRKFJAYqlVbd4WoZnsccxthYTweekz
D/dZcHBs6Fb8WtM2DEfE4Q34kvFBHQR5eCs74E1Lno/rhsq18xHQhGfgRtNIpx6B
CFXwrmZHsJCRWIKIAtZT7vJCK9Ym7t2eXPV2w35QXEjOOn9L2oJnXK8XUjOCadAp
0mqdRAA6isATHu2SJSgypeRTws+tBImKVZnB4UfEnOIjgmUyH8vI5iYKKdT8SqNP
SR9qn6IGxtsiWcLtBNL9H3P8r+S/FZpyuz7OAzxdyYFko8xDlzaChSAs3mOrRn0D
w/maafnW7e2t8YYtL6L8NZFClv846CRfq/IXb2RcBvYsXwjrD1KAOE/1/vbNZCy4
8GRR/njVPgjwNU0fdoJwhWx/CkehqhTsvF6LWnxZPV/Tw+1EsD2YGclKvsfTfCRD
g5w8mXwrE+W7pneKCvR1o/45LbIdz5NUs2g0iia8cuV4UTTen7azgDlozMKkz/8h
ue/lK1mc8Ri38URJnhoHCSvooxp21X+0YqmHGyIsQFqrLZMyYOv/Jg16l2gVCSog
q5PWXHc9lX59W1EzHENxy3b60l5pp3FQZ9yG5mWcJfiz+uuzfirtXTi3rq/CTX2t
SDbRcmAUjQ3dqnsRbwNp2ZqIQb7Sd6EiIuhMiHDKNi3OXdbrbBwbxH79UtCX+e7d
ixfAbB8+PzxlMqu7Jpl6xxkjBkywX+CUftEV88nC2s8Uy3kWuHjhMz5kxnDBX4eZ
Y+OCl61ctRtrsHZdDFbRKWph2ETj6uUXJjsvvAu1CGL1COBiFeACfaESbOWsYwWk
ttHoVK5ZGsEUw6pP9cTDgtVjt/CuWDH8J3CGCQWRhHtk/yh67wI+zF212frp/EzX
i/td47mKST/ojd0xsksW7EXElp5TkH6xCDePCoD3dqUQZnaA69Si+PqAUBlYi4IE
MLGjj81Jn0fTZdpQJZIyqcS2jf0YBGOpGsaIdU10e3bZFMCyRFEPCTwwyX0OpD54
h34f8UkuD+PBZ6HZQYI40vaqFBXEzMb0mcgx+3WvzTsic9IFm6xZEViVN7cPXfVv
DVeCFBY4VZ4REUx84Y+Sn7FdU8NExw8ztkbsxCJt1G6K351Le0XmTs3OPfjhucm6
eR7eP9nVA+/WsyzvOsqETYfmZksVmk7LKMld4r3wuGodR/9kEOPfvfP94XoI2gT3
2OBzA1vLqQY9iMMJqXMnyHTvQrkg87e3Y/u5EWFuW9LQ9HoD63Z54HSu1xUHf4kF
MejsVGBOjuX7NJkHJrIwPZVwEviIvEJcLQrP82kpwCedpBftRqinmpEoWyenucHc
hxZw9GpbNg54+lronue0pgXBF/3t7uTJK/zxED4qwGzV3NOpG58d8NwFSm1S+7mc
kIwtJIKsgI9fLxaFZcw03xbfUsSdfXUU43N4Qu5FAyniPauYAgE1rBKVyhhOC+RB
Jx483i21qJD914SKmPN5303/MG6FJjZW2cYgXFAHV0UD1W9x+PRe4C0P/27dFSW2
d8iRExqbiSGdzu5FME4sjJMRleVmG55QT0v/JIhvrJO7nfIBGBlJ3lh/0fOywYSM
0CF2/6vU0BLSrGqiJh6xKAAAjx+PAfvse8qt2/xqhaaqMSQJm/d0EP4uyCoGZaH8
8DnwdTasH2hvD+LIwRqMvDBiNz2zwmkVowDAsBlrB3XL9+UZqJx7EWrajYviQEO6
SZKHwF/7ryikg+YJAj8QDlfoMjgzRwb9PTnLkA1OeeRmMLe0NHq9205WQRUNwJEE
EQ6dbEl7iHbBxdzyk4JglJ9UtUcQ0BAcI7scDcbguqIUhrsk1+tZP09kSrpoDI92
w46zafDRC7jaMG8fGbaCfnG4RmimE/vsZrNWrtaJfTAOAWiRcG/4lGfgyPZLr3KX
7QW5Ns4CXE37ZqUTzbiRBIRXNlanjWIDpkQBNHP8ZG2Jn4CDHQupYbX40z5uAAMz
o/XJCZP18sfZyONYCQJUFRMpQqQ/0B0iWHLkYKALXsY+FyWuuJ9Qjv5UlEw0GKI0
xEgwScVowQBeXHahYFUh44epMMhp5ZKSY47nBoL607YZj6QR3ApbQfJQtmN390Dw
h9N/FVJzu7WHNfAJOQ6GNxkQOTl9NbKxKc13ORu4mO54mzUnQJL+q4lVddG8G6dP
rJpJI9trqP6k/aFOabjo4OCNtVWW4C+56tmMe1t4Wz/BqSwABG8JjO4PIXSD3XAQ
De9X3ork1VzwYCoo/laKEX8F/99SU593/ckYg5mqZ5wIujU8btGg9Yxe7uIYVNwK
MsrkvfSQQWQoIYAhQKlNjQtfe2AOGmJl0o8XM0zzZeyiVCpnqaAC4uDzNsIixub4
xfkd6NWTf0/ak2f4to9AxHg91yLMJjo3I1ocH1/Bt1//NAXpPOAE3NYX18l3z2Fn
k4mBUCF/5OakKKeWMK5MCk+YRKPjNDKF60LpOk9Tw3oZOFzd7TQMqEiJ0AnhUf0J
NvppQdGshrzIfXR6+EqFCqp7y5FYxEYpro2/cElhs3eAc/UnCqu29Qjgx1PjmRDu
MEubtuJokq6SYVq/x8g4nj9qftraa34Q2crtp+EOmKx5jXfsgxC3Ulbdade/LzK4
iH+qm4oLItFiMG/aV1gWm9m2mbRP/Tz3Q10LLOlBly2euG5LQ8bPljS9DdJl1RDk
DzGN3wljOL6JAF+byhS2vlOMH0bv5WegSiVAax2iE3PkSvOQf5LLfHBLU9DiN2Ks
25SCkH63/2mpNV4HA+hZakn+ZshU/M241opufqbKB4h2z9s0Rs/zDcvjdkzRT8Um
c2GMaR6FXA6eYN4jrkQFDXjstPzQAYh2y1UnUpgcP5V8jemb2Wys+1jsq1YyGwqD
n7UA+9DaRd9sDjCbEvVIrzUYQU9cbmlkOS5a3ztkav2P2EziTDbX6f+M30kSPiy5
+D+dWKrhOIc/n+EfoxgqjRuhOjRuTDhpqLm2RLySATZYeO4gzx5fdLCbKUZOJS/V
dSaXtTqInKFalKSlwkEkv9EFwezCQc8XXxbDMp7MU10th/L6IfbABGfuIPxaiMIr
0y12Ur16neIH4I7ufdjUiLpkNNc5WruN1XEXuLVAYyV30p1vbnelzrfNdnPN/Gi4
FKftnGPZ9ZLLBkI6Sj1CAyyPP4AtrvhHGHg9R/T+Y9oU8fnFDiqkH9GKyJq41FOU
IDzDtO7Qg+7d4R90vVE1yqkAMmxBa+InhkFwDyK2avDD0NnOZT6MPYQxZjg2C5tr
kN9txvEOsz6tDgoxvR0cQEN5PPiSXi16unIHD5MtMAi2auyNquhVT9W9FD/bX6aa
8NGSf3m2+TyNBZHOcji4Wp+iB1Yh0rB9GvzocSX5PVu8VkbK3rxLyoddwC91IaxR
v7JhagWvdOEqKxlsB/RbZv56Z7ZBgvOnLuCDH9d/4Y8WC4mrGTMB1DKVmx0Ey9qd
JkeKeqHe4ESjpw0g6WPjaupvHwL45Kc4fuz4T0g8LLm+Fi94gYjxHb4f4pODLz15
qu7kM3AVYe9LFadDPZe6KZC5x7XKNecS6oWojWm8v6Bt6tOac3uykCV46X9jxWrT
1uDPB+yaeqPiHoYSAOdbH1s0ehgiCdhtSnlgoShEQtr5tifnyIqk7Fabg0+kBftb
pru/oUtbbCLRKArHhou/m/7E84In4dfBZXvoZfBnOps1kSM0UiRppqSUfZOnrWey
thJRcYs1KgdKW7Fhu6k9/9i4bttlZNbkDpWFzbNRamB4DRJRC8ev2fsFGh9jzWLK
s6evNEzvzSyNRX++055xrFYnirMGP8DGfr2IMHkr4QqsoO+WMkg3W8hb/uivGPDQ
Xc43Q+AG4Tdbn4QhJwahuIKA0HBk5Et7c55O2oL0GhA7IUJf4+CtPIszSVRwvZiL
R+Pg9ZPvoC6RfPTClcjVLob2sGJe5uHqBWCd/JT17gGM+HI/+fUMxYuVEEQuC9eC
tvlqnamNglOA8m5FDSN8nZURZxICM1K5Pm41kyum04da9IdpnilQO98lsZ1kvYQS
e9XtPqUhxo6YcR4Daheejl0vLVW/teVu15Wk3IXPvURNeEAPDsdni9rGUbMOXHNw
mc24zFgVtlEJzG9sz6dq/J5pvAZAnw9Ok8PQ+cfJI3jmFaD5A6CYKmKJ+Y/GhKfB
zlqKsvgQLRxPtPOOYXnHIzFxQuPvbGB/IOwQs/sBVoNcHrbpVnT3TR9Z+Gz06Wpf
ag7tUO0ADOQ8Ow7fnxkFiEDWmm0TDlNZxm0LblrVa3VtDpnXfpJ+HmqDH9q0IuX2
UDne4VFnWXE6q83RXK9GjENv9nmY5zuUazK76te0YiKrNuZc+OL9SDfTXtBsF7Qp
gljk8rosAqSl5RiZPNf1mHVy+eUEZiMZyzJA/EORNqp2RVHxNDSIzHmomZr2g3nA
rXr3kNJ/CpnDJhrM2rd4a+NwFnCjroNEO6rpULR+z/hInJuq702n/mT7c+uI9dBM
prm+1axTawbn7GM8sUk4/fPR2Iq+u6Y5mDH+KoSGXrsK9xrVoatsDMDflQzv7SEf
buLYHLjX2oz4ItzQG40PwocyYPzfIcIIi+O/iKYgN+sSHajczaWDCQJQc+BYwxaD
FoY8/kjt86pDz7vfdNrslswoWQnn9I7gZGCWk9Q2qzOrwysJhLeup9iADJOnIk25
8oI/HFq4U7l1eGFGZi/lcA9GMpprEKbzdLwlrHokQgmBGrD16d7xFx8Ktxz5VFaQ
kIaseXxhqeU/w69Y2/ZC17sCpKpL6X5TPgDqugFP+RT5Q2BqtcUkTbSUdVjfx31A
F4j44BbMjmQbaYqLufRHal2s/tkNDtjpwB+DKDpqEFZfIcgBr2XSvyXxXYYvCgtx
piyuAV+QPvM1SjHCfEpJ3Fx9wtx+3PBbTpv57DAoD8JRhHK4JykhwPIuy8QtvejZ
0X+GZOYO2heWJe6nj2iEGFRWonreT9SnXgebyW3Q1YcWPAW2yfez+Bheg44NrITt
ZPhwR17P5IOlijZ8G6qcwtdb46ovhjE+ol8VMfWRgd7dGWWjHt/aemeWkt3TmsmU
TUjzWVB6rePnNet1BuF2sCg+VpbSVuidcMAbg5Zlc489r43l3vZcg4DojfZNBPJU
VZ3DIMka3HxgZDuEG/IW5VDF84Im8CNja6QlGHwqkRq0Q/8wg9B5XefN1ZvnfU7i
vDs7KK+ig025nVsUIXWJGWVGHPp1qxUrhPU25DwvCkmk7WEEwHnQDf7JSqt2UDEs
PaX93x0xg5doiupmmTgxYAEXoIhd8WU9gF2ugq2+7tK/sbh5aKfvuWfxZK1M5RPm
CYo3BVRvJSeUNf8e/cn17ZaLOTXE42r/EKnsmUZMcxTzaXTHxqM1MOYqPUAaXa7C
DtD6AfDRi6jssHfaf3fYo6hZqulR4VxdLtzk/+WABmzTHZdBbJCHRgwEtm2EaoOx
v9hPDh4DLc4Y7wRNaqOCIgQ+l37+IN4LpLNHuq2ZSRVX+DLf/D0+HeWoGTKOBa8M
echoLtPgoc+VRPYPjQE81ftu0VqDDJm6toP7zdLgWTYadTCsPzStgqOg3Od8Nwb4
YZX6IxfVF5PGjQzNceqViLYL7ysKkW6bbBrY7vk7uOVP0bWZA8fnxFkNcuG0LS0a
DUEtUSlAP9biqz1/jMJFS5neEea7o8W7topmZoMeTnzK6Oow613HlF94VFGbUbmL
PW7xcaGgjO1LPtqY1UuNYOedASG2fkXjNq1OCWveZQ9BPI5y5Q5/aHcAi4PSHz0b
L6JSfyIB4fEjfG/Npov+47UuJ/a65ASQp1d+dnMHZxsXu04SJi21TtpoQFiQXKPU
B4sdf1UF9EShq35Ree6GHwqypITC9klrxEAYcRjWNcDHN6OnugzIlhpQIPm0/SEC
eQlhrQiJV2Mia/9ElWiXZEmNCczWuvbbCyfLEClwkoGHRUmFOjoKy0NC0KJbkOcs
k4VfbSh/MwY0GXLUk3YgI9dAA0LhVtsbjB/LSF6o6hpIPI6tnX2wzLkX34ql2M1k
DXeggWFSGtKhDozl2Gyj5zsMzQkEddzS7msnd0+QlQ613aypXupAxiy4l1OOnWEB
xR6MpmpdNPYqrT3BwAsEAqaolyl2UhClTLSqKGRDeMRQsC5iR7uaOcXG2TTiGlOA
j6mCNDxISlFHfqT3515Rf+3AUD1BHltfSCeh7LrfFM9RHS1cp3TUBIcCblQEguOf
v/6I1OwuNPt2/hrC8M1J7uC/4lt4CIjqQtGMSmddxz69KZJBS5HesySfHOBy0zou
uismk3TqGoF5bzsofLmwwBhqc4yvb/CIx00UOlc4iVM2VdJ6+blFV8QPhqkMp0Rc
ZpEHcAsuha/wNnnt1lvWKR/m11wmKG/F5upV727oT1wUsYIpyi4Iqa38wL+C89PZ
41ntD4D5KG1Nx1iZHXK6h+mK6s69M949p0p6SU70Em2jcTdny/by3j/Ltc9vGOWC
rGA/Fx2u4RMX2cMUPRHXq4hs5wTd214QIo+uK3SOqFznEM7vPGfq4AmZ7dMUpMuW
QePrCQz6v1xMXeNqkIPvf2I5VJ9018Ti10jJaioA8sxxC+jcnOLPT8kh0y+0Q/kh
xOs9QyLT8neCJSYLMBQkF3S9WAFXn7nCK0O88U0DPtD7KfwCHvrCOgVx9b7OlF7j
SM7K1/F+ZKO9sWkJOFozfuI/c7ertAOKoPT9iULvoRijKKcQtCJsDElsHwSCsa1f
ZrQ94h55G+RYOX0vvUnJgbeE9KlUCcHiiRRywMhffgUv8o7hc+au5YksGWLZ5pns
rXKtN+dkHvCvd86G2/BXfhxMXWgVk+U4K30PHoFlrMSTQertQ2ourq79LEI5gpit
Pvr7uofYPt1HSG3o7byVfmPcKrRuRwvRlvNRg1zrhL6bMAIeWtEEa1Yb1ghLfKzd
jsYFZBpYmFZESrK818SMbMU5SQjh6N1Dtq9uYn/0EEFSkOAxznCq3wPXdXbAbGON
XcZWZVIYShtWoXJbi5RsRZIiwQhIDJtnml3LFvB2JC2AQRIVnC3+/B6J2TPHMnQd
naHL9cMKWxQiXdwFnfmc2jp5Ykb5ERrk1JkM1Jrm0atlor4CgcudwvTbLQxGYVSQ
MZkZBqtHhngwMzXf02osI5H79RcNheRaSUztRKBcnMtrRxq5o8uZ7uBmDCew1uXy
8Wv2hLMsNLRrvgkX3N7NBXoob2shdgtOS+5slrdK33Jh6+9r4Y6wyRdcfO7zmI0C
YhbyraxYVPjJJy1NAdbMejPUbDNy+64FKQGtgyxAw6TR6o5PCl3P6t+bZj+ns+9s
83yAN99CosCqQEOoplM7kLWj9ZDchJSlSK4KaeOCCkDvbBBFPRED5QQm7iQICdEh
xoG1fpuozOOy89hBMaWHJG4PbdjMQAFBl7y0pDQSIi9tl7Y918cO0pDW1Usjj+AI
xuvSDAL6tzdu/dUOzCSnm8/ivnmrVdrIxltkGMU9GS5FpZHNWBUTlHqhDlQBb5UA
yjV7Jexc038EUpRDwjQVernPAteKoFWhMDi4cAwiNev++XU4cIiF6PjtCpR9Tjmk
jzUuLq9ncVuoK5wCakyfKIksxDaO3/0vGxzW3hxwfhziwaTOiFzZVL68g58l90ur
Z8ec0ascTA7BLTo/XBFGoiqORuDEh2CQPDXM0v5ocA6NK5kaumtctWJGqmCjHfO0
HzXyWTuXB8LPXBix5RER4pAQ+I4JZYP9ropCH+Yvwo+N+t+SA1eqOA9Rsid6CiBH
YsmrHCd+i3Edi42riMMHNQ5w5/CRZ+hzDmHQlM4BRXRXYlG6pvtq7gAubXmYXCYK
QGfKt+6SX9PmjhtWmHQF/B8qDIQ0oPpLKOC2txRKHT9Srm3GFSVF1WSOeAarAmYW
+Xono+LvIdWBZpd0Dcmor9Amhujh8OYgI4saLbEMByd81aWXAsU1TOHdLaUEsQ8y
dVzz+850+8K/pm9+IybflEgiWYp/girg4M7K0FzU8PfwszHnzc8SWemkPFaEmb8S
LfWiy9J/HTr6tkgRxGxpCUXsCPcwH68t/29pKCX5FneArSNby2cAFOxDrNop96NV
qx8KTsExYuZiSkkSq2SEBzcRe/GIjcCMZbjsuo00NYmV0a4f++tP7QiaWeVhgz1s
HdYR8ZrTvOuSRXoCyE5XoGhy1Dk1tXP7R/3w/zOwKsclfmZJtayBFk0N9oY2cv/r
R/R1H15O1Enl73cQRQ4Hi4fHfITreNME7smpMSP0pYzTgftgZFeQc/Oq7Ro+cc6V
pKwed176RAdgvOJFGQocvOBGDGw+DAb3JwuRHFMUMMpK790SZEoAv+gvonoU9rNb
Xv3aIeB1piwKSmI1Etox4/gHLDGp+kQ6AmQ1I1G9cil7RNQesKbGd5Th2IlBNq9z
2FY+WsOg3A174r+E6Qxxhh5VcHfI1oO/tX1Wbl7ghyx5vNuPEPurub+Ao4PvXAPD
0gy/lGr2jxlQ5mkE2yIdmzzsdoygQ2jO9aPMM95o6py/nGe75YZJMCSQgD2xEd24
GM5Zr5iGHPzRP2GFyDxemUwKh2Oka16kLrup+qxTU6HX9eLCtJAvFUFpEAQ7wNtI
mOu0d3hCPrRW+5O87flhYrJ5mW4gH7XoQ4RMAlXamHwz9Xiso8auHCXJWVT/8ZZv
/5Lu41XZY3ilXhH1i+A6PrbcEeiGdoL/mV4nTtNRd88XoOcESWEieq7tu/PuORGX
uzZEB7DPLJ2ykFW2cK0H9X2b69Dw88EynUrUE+yKnabtWQGuRlzq8upOJ8ic8cYa
GWONrAgSkpwROfSUiHQJ3/MfsM96OTiTSpX6n9Aonybt9hEnePzGPhY+RcqConwr
nQvwKACOOjXAxCs4dPEJEZGS3BxS/L22eH6igJgB48OuPXXtpuGrBybrKQ4m/paH
qO3ZWCZXstrrB6d2V0ruYzlrGWj8cvhf+Brio2K85q4jqzBnUgNqdU5RTIi8igUh
YwuVdIlxdXxv5mzJSYNWeTONZeWKHv1ARa+CbvhIlQkx+EWMiQcEYiN29sIGp/0P
6QTrlhm6TR3h94Lcwd7z22HvQKCqY6Qb2pBUDN78DdAWUMzJg26KLpBf4E/C12rc
DWJS5/9o4S/eR9ICwH+Abg2dUismSniLg3iewfb4s/o3k5K+tsAAEaZ7vHKiwHu6
fptw++OwAkbmkdldyplD7YL9Zx3yNDOjMsEiUHQVcUMSHkazQ9gaUk/ZcXJailet
3KIGsDaSY58xZJNDC855Y3bwqR4z0HTgMWij3tEgIIVItyvg13UwLacFF7qViBiW
V6nPHsaFDFDV3WNQxScj9uQC/yMvdpaeeQFnBIWaM1HRvX45sCjk/GBdtxPqV3yk
jrFjctNg9LWl+RDzM5Qw7AHsSXQtgb031iitl//5hHoDMefP7jdr+998Z6lFPB6/
4uDH0DUKUYJlGZ53NgdebOEAU0lhqwEDDHSm90vTjvg8RhA4d77cK/LNbdEdH5Hd
ULOQNiZpfWA/fSU4KSPtsSBHXeVmkMpiuqLb9+hcj9MZosh5cBjwm66+Id+Vaaj2
XdjaLqh6dCfBTte51eCSffic34pJdvJbAFhlMa/TCG6aumlU3qryOIigwTgMEBYG
4e/bz48eJD8qOaMMGHZqGrwMG7DTxTpC7MMi23vy+62xG+N1bFYg0arYxIzddYka
8HCLk7G2QSQc9fVr4nBjSYRF24VG9wpC0bPe7cUZz+5bexfqI+6HZUYOT4uDRuar
gBgi8TZ6Rd2RUSRGcZTWKP4GPLYmlLLwq4nrpqZI4A53eEriXEYSE2tBaH66jFKE
VYErG6sTcnc164s05QCXYoU7yK8QJkGGzy+ZkfS4XjN3dvnoU9t8yINau91rg4no
IO03GMG7oWf1O1ZmWahe5wU0NxX3dCXFshiveaUpXQX3COWlxCaHFBzSCIOfVh+o
mHWW3Drc3X4iiW/9TeydX7tJFZky3oKgI7DeYBD95OcHZGtXfK5BZuOqDQSuya7o
+oC+/kwqz0CoAOgrtEPyxuz1uxl26QZluZKesEvs4L7FrpCcWlSvDgM3t8FRie5n
mlv+rxttPupBMvVPABUsvFEj7NbostgmVy4BfA6cWRbUkTXaoD3cC+V6511mvh/+
xA5OT0wep35FT3pMLXQtIShgobRhW/gx33SFuivtDkzEnroeAU6xKYc+7dxcxYHe
trSCq6RPc+vhuclsv1gX4OPu7LKeOoUCP+Dk3BBDmgGo8sKyDc+/HQVATyPpjbTk
XGpvXnFOWlIejJjqr3vLiKeeqQ0sHAQm8CPsjRPCbDfmh8NMp3tPnXQdVkontNhg
aUtW5M1gjcnGcg/3VaZoiI4Qw57XA68nYVg5KVvonvJdltkuU6Zgn1ymcJbp24XC
blT8fBF0Jt6skKRMy8csAG7R0tFL5S6QXArSdkX1e0oLO/vmA11GbdhyCcSkMVpz
kUOQEZCZZzV1BsVdagZd0dKlfc7SocpQ/2CGXM/IPBqPKTz13Cyh/QCQaKrqfVev
wcmOXssjI/AFQMlSN5piQU/8tVLoKHtwNfDXOGeJG6EFevorBzgPGXXg1fPCtF3w
L3FuMV+9BlRhprD59omXfL9RuQNGOherGwg8zLn/c8JbvSQsAAkeIoAmB4hBaJ84
mskTqDVBRSVwNpCxM6kciBdM1hAIUMDkv6Ekb65++n3LwRSrKi1TBGbNZ05FpseQ
Had7fk4AVITcySzloGeIGcuHQ64SO+5Z2NzCKk0JlAxkxmqkaihnmHXXx6HBIoOq
YjMgP6fYt61HLGVbvK6wXwUH6lG5gYXo/9y68ZUoiSMPKkb4eRnN2KcInLDPegFS
8xfsE007FYbnsM1LqnO7X3qiC3mny573yOYUen1FdNiAcNeMMNYRo0RJGkFLeIMP
F56OSRMO3P7n/S67cOyr2/xxAxgqJ+ihri2cR9Wwen3vBQtsui9vzSsCfgkicyvY
xXsuX7GYX03JztfR71AYV/yYqGTJrHtHJA2CRCMJOs2WTX9CvCelOiGR1ZcVyKiF
+tMNyiLafVYCBi0JGqminxirfdVN1AprmCOtW9EObSfWC3E6RYYk53w5xz2dSJMn
j4LQ5IKoy+Cc/nOsXnWGwguuPn8Ef27ZjUmTucBFVqO8SCLvIeMi2eHxaFWA2wQi
azz5SChRVjdNhqt2CdHaV5HhrsX0HFJyTPlfWxW3rCxSjTEjw0uWioLnoqgiU+rp
ykdrDvGBfeSj7yec/NFAWfBXWS+IUE1PzT1i42yiUEAXOO37urM08w/wIaSgoQ9h
0O4nNVZgeAoVO4St6UTT1p5QJ9TF9lIgz3xl9/XTxjiAWERcC5TNCnimmLqR0hir
VyUqyx5vIF9MU4h6u/7b9bpvybNSvr+z1ejKOZC05lAUA8/YJJBO7Rfj7uYpWPa4
YJlpbmVamsoxIvixIr50bfp78mCqUYXK28OaFhVaCoUz76ZhSf5HNnoHbiBcl9Pf
0J6nJlyS0wRAtJcFIx3eC/A6upxtX0SIc51Cm98Uczq8Yl1cXteWqswt2GLbYHWn
6Xo+eY9qnLWuH7uBWA+x9j6/zF3FO+5LoCUnpy6527skMvwyRAZes7T8tu6P0d+X
sVI/yViREwc7dghEWzo4QLhFx02tXEJVTFdIPhl++lkCxx1UUwYDPfCDHaFFSG48
stX5uACUUtgVAnd+60N5prjSUh/re39mQPr16bZvDtp5tCIWbNZbQJRE1p4J+iqk
aNe7FEeS56XF7EDVXy/KFiVpRo1AI++4T1WOjQ8bCKrMglssgg9g8hYVz7qIY8hT
Py+rXERpysr+5WZaUkclSANyCkaFTDp3ojlk3ujXDp7YXcu1W8AmgjZyYFLnHwoj
zaeOZq1dpZf/IssYs9aWn5BPXQ7cX2N5XRH4Bqt5k1S6rzS5c95k5Fz8qdu5wFfL
0vay+DLXbFet4exT/Xx4wda90gAhHfGfT3mVlFWMUwsVeaD7mul2JXDoxEGD3+5b
ztm9kQ+Kj/aUxi6MRjhtOsJ+tYuAQBIxyOn4yFMYAqkQFohnkhydSkgB3ZLwWRgU
2j2RdgjJ2hXr8+EEnVvHYQ6ntDYhsIHYflAmUD3nvkPNrPtA0TfajTYzn1os85ow
oD22YYW9tzaYrAxnj0g3CHcbhPdkHr2g4XFwXBpiJcTMNjEauYcQjtyAk9mnZ231
aX6MYgdLfbchU/8u+Ua061SCwMmxWfHoBMNV5XdZ5Xm70/vtGQItYZjYYH+LnOqV
v2pFDKOSXYd4V5cmqFGM87x1QLoBHIu8uWtVn924I6DMfdjZBfH6P6+dnVMF/Ne5
oee8yjgubp+CmTXRurAhZBg9nZVcKs0NDdqg5DvXWR7RUvWpx7oIk5uOSYO13xbO
FwwIzXjvIhwbyCJ/gVTHG5pjocihLyUeu7qJBAkfiEuzB4xZC5JqgsuLF8YtO88q
vKCSu9i3Xvv7QdVhFo5GPY0qq5gcI3oAcEArlvH7IkFu1vJ0HxR0kiPTKm6DHn9g
3Gm8gbbxZmmt1MpSzM/JgLNkpc96lPyce/YliD5ey/58NHGt+hLYcIwFruusZGHG
QIhEkEayd7HuzyrHnVoOUHnYUcwf0xkpL6FfQn8uDe8J2dH38eij7Wm68+RJUTi3
S0k+kGY1gBXt17iH8UUXkbb+fIgDYpxVXoEQr0WhCsYuogoiMlJk64cXB0CQRXcH
Ja+1KrdPbsLkBTYj0nNSKbIsXyM9Y1zMtsAUcpEWQp7j1njZFDn3bycdZfxkv/+C
gH5OnUYBCqSkWUZjTxJBNn/V5n+TACRjHKSEgdRDCN0jjsRp/Ldc7zhyKR61+ACW
tsw6wgJHLUjEUqOxDUtNmYzY9dA1M38Nm80nLSjXxEfQAK83fvIwi3hrYEskzwW7
B0OczFG2+MDAb1luw3IpScP1rpVHSj69zRsupCI26YJcgCrtKJ+Xp6HJzOEZtWgw
2xYJpcWqs4abaIhRfISnDaZWzflCWMbCoeo/XAXdAWiSOrPGzbb7b0VgN+3W/G3O
W75P3SxwYzosN7sAwyLyMfAjbKmbDArdEEKI3ZGb2xRhhEl15Bs5m8V+S2MKSNs2
S4elwDAWVshJ3yuNS12YhNV6IGDB4VPCHOI0V/NZj0umZlf7VENjPq6TmJAwH3tH
3niOqrSbaXo/ieZRkpj1EBmeJAm95Bej/j7dBaD67v2J+x0OUcFMMi3+39xNRWmm
8DB2+y0zhXltXwdpTft7kdJYAks3YuKMHHGNKzEwZrEbKiqDjP9XPGVU1YtSgBet
BXgJygpDVfKGztzRj7LNFxebLNxLVMwmsF/JX/48CngXn4uE/tOYQGeGzbxvWODc
JLcEXmkKhxbaXVT5F+zQ8OKi9WK/7GEunU7L/dZEitkAlZfMtrKrBPIrT805YxoW
ZnsZ7ONx4OmMz7oQ1lway1JmdQLpm6uK0RO2hbtJTMya9UK4ziGnbijk8eLjJCsV
sI+2+D5Wrk+d1Q7H57hrHqJQ241eqhT4hdhjjYpOC+WnItP1YUVSa2EtW8pelImF
oe9QUrYXyYnhFiXe4LfugPSjp27Ysz4O/y3wW6gZqRFQ6O42z0k/jwZeinci10nU
i3+Rknr5+ob/B4xG99xn5BxkdeMOS8CCReNxC0wLqDdJba3mI84SGOfZmZBfKZu9
AxSNKFMR2zzbUr8pIO8GxfiSkso+ZD2U1lGvkJmKwMdHVZ06dte5z3jz7xkMiuib
PF/WXcIOyWoT66BhKkJmITZqOm0Vgu/ITAnpoUEr8MKRLsBYHeZO1p050agN/lpW
IJdqAofHuuUM4huJbUhBZPKZZBKq4LApAbRPfz77ldEGc2JbDsM+GTN3BBBtZt8L
S48fhKu7bPGjd6iKVZqhTt28nqRndaMq0v+JD5EigrjFJtaJXHfXZlzNGAPEypFG
e125ZqdCMURYpfl4qhsdphyZkHV+bIsxopXNYqUhlPdVHDvquTumc8pezBUOwdB7
GaKnrWQpwYdfaLPj+n/ge4l9Aa9k8hRZ711MphRhLoB8gGE5z3JY1VocjdaSEb3I
AgAjfOQZ5vHpsey3TPtm0vyF/25Bi87J6FD04hyUirlSFF62ekEzCoRqAcpyZBAg
lRcn5iSKhp++7isDbPv7602OgQufzG+pf8DTsKE+lcYYuG0B1/5tPkH4Bh70cy5G
l9sf8plGzTVwCqrmEN3ESaTp8TXEPekqPw1CIb7H82IpJnouEI0jkIHRt1+9lsBW
8G/WPx03PNuCs1t3c2pNCd6b6rJPgeL1ZWUe+gU2rl8Gqx5J/fTi1o/kVCQBscZ9
LJKV4YorybiAJm4pzTKaCVjShxOK75alS7zEcmgJjUGw8JdscefUQr3csnW32d4E
QX/wzUnmMv8gAOUVSTTSJqvw2dDy3Ndizjj2TbONI7c7xGrKajqEm+562I0hZzs/
mI0bg10WZw9GnnsIFcD9IcoRFCuGadlFBW+sDU4kdNkuiNLFXiK0L1caBjPUBSGf
7c33UL9daw1kvrt8OI4DW1j7CKVkSAITWFByeAgCPm45K1tNMHggLR+3jxKfOZLL
YI2h0l4/UUeCpZ+VgDRffRtc9yDwZJeUaWByqpM1SuS8UwqOUCbcvyI6OPqwGTVf
M9OMJodtQki2EgEXJw8IQg6Xt0RoVtrJIPGnJ4FkvLbnCr2u68KVjp9No1toCUYi
GjeN9qA/Fda3sTR4Hhc7vrOsSbAZCJwvGS5g6mjMccck0lEK37RYt4Z1zUWMa/fM
LZyJ7DcM0dGHg/Bs5K2dkuKTBtij9IFhAOJ70HeNXSz1JcUv/HMjV3DfY05+lroi
OeVAqQdFnw/Jrb/Er0clHG2flyPlYPQOwBAre26CxNYhNNfSPbLlj/fEanqVmXqr
cK0JuMzsTkiurVYI7z2FWHf9QVdz6PjCFXhZ7oZWrQ5xBj3rd03CzxMGsUyCDezR
6RjhEnq3F57/8EtVOq7W9edtjk6n2QbMowcPBEZCqpji1Jmo1oISsVbeOhtmEwmY
stsdDdJkbl6nkQy4c+9h5LcBEjnTJ12n3a71oxFLEKUWbi00AwoG7CtSRqJGbUdI
aXk2st8p0DQyaEgzLZ2wSrdiApq49tlB/Emxv4xhLrSq+lAAvEVaBVz0fkPLYHfG
6VYQZzFsDEBEUtL0dV4rkc4cSWsoZEQxjPAA6Gyk0oLOkyLSUXyziRY2vdywTETa
zuFFtHFsgM3UPuK/4KrgUWyFhPRN8VpLotruykTnxprML7pUqywZTiW/jQfmTd2N
pyQmYTsUyjVPmggY/YFhFg7X8F2If9k8DHrGldColmO8E0v7+UhzQedtDyZIRbt6
2vG0lhA9MqR7TO/lBEL8yqLp/fclifFM0SFW0aZ8mkAgUOMIchzocPvLArwDLH03
j69olweQTaXjT4PwD7yVdiLTc39Sc2nbdtLmOx+D2wKLL0Whw5V88P7ITbzokI6J
mb8ufHIC5Mq0x6YinRFpIe89hILXsSJtX1+K+SqYpqSm5pBp8PSD89pJDUshJyRG
F+vTFC8ner9O9dRi/IKzW9Q6OwpYAzoCIe8N9tthowTSXDOte8h2yLEN5AYRBJ0b
OQum3PBFgbDjirC03SjgMfJ0jTRC2o235MeWzGoZyQzUlPDgx3w49k0ZZ/O+BH85
z6OZojEdY/stbkRB3bxuI/sr2NMLnezcA5DfprR+Z0/FKftCSVJCJkmmYeZQ5SI+
RVakLWUXFiLuWJ3xB6/bEcK54x9u/c5qIrB2rhS6FNvN7hYevBZ9hGpRs9JHN1Y9
JlogyJdfe1NlNEuxvdfqY7MKxlVo3XbgBDLX2MIn0qJx+KCFwMQMKrpcBm8CrzLy
3RL0MX2ONnmuxC1ybUsMvkxcX6StMihl0XChioiYGS7H2nLk0nRZ+ZiXopsHpu9m
25DteDWE4K7P2qYeAegqVAw0FIRyl58lwnMttp5tji81z4OYm1QVxp1d6/xALw+C
khyXUktQbGqBDJO/lnEzwEH4D2V5D1jVbNgsRsUE/DUG72vxVEFVUExJibdK/GoS
NU/dF/GB6FBpthotErq0iq5KUaHTnCYN58fL66I9LwEK1FRHoE2NEPAhwXLWTfnn
k13aERFPeIgyuaO+2AngKsqcEsq1YV81jD5p8HqBdnToWWq24npb1TiglKdnrseL
U0OOFGilIh2A4gBcwghYL4ybWgX1D6JgLGBZd7kZFOnKuEgzNL5lJOrYjDbta+se
yNsx70vvmWoz8lBD9PmwM5q+9NCF8GsOFl+0blczvG5iFzDIsmW5uTFb0wnNRKFt
DSzy9PASqy7ySuFm3TYpRXk/0a63epu10zx0kRmEdL0xbl4G32EaAJ80R0PrPQhS
4LNfkmTyUv4Iu4mhXdFpmkuTNm+UfJ5rfR81AbB1U3Z7r6v+ldlr9m2tAD/36zvr
cIIQzzYuqIut9JtVzvjoud2hiMFnmqQpTB+g4q36aGxUpOkJe3j8AIHTMTWNPIqU
/DwbGRrNHjhATkAeRLIKg3XAJi4Bi8pcCyKbpqHnyhGHM2TmOjfx/OW+Yp8nLBdT
DvuqL4YCZ/ge/sqDPuRcF1egzkBElUX0fRjhT6xdCA+QuI/Ng+TYwLnpuUcemC4C
I0xWHr9oNfIjELfppj7EE7LTanQkM6xQxcMXwFT3RMdfeoDX4AOJD2q133tw6ygZ
JVTVfdTsfZhztUwHr2EIFO8JpW9CAcXl4dVbB6k2aYtA9dxVY2poii0Mg87JMCjd
M+ZFo8l0iDcUibFWJMud5WGksqOE828MzvhlVVgOSrfn58VU9MOI/B7tC1S/bkkP
blol7yNRuYurayc1zsxWDwyMaSSh6HNbcJ7flbLbBzK5vwc3cxZtjm9q2bzqk9b0
58lMHDnhN2PyyGpQW41b4oNyQR4V9O12RmH5wjFQtrVyFHnm0Fn+bw/KHttYAMRJ
UX7CUucTawLr0CheJ6skEWd6xY4ilYKZRPoJrBknL1fnA1MeCu7MPQRWf58nNJmY
Fl3wqduXiMsWrfdvhsdLVU6MIvSkNObmGE9AeGax1XziwVAKp/wjBF+SUFeEnHc/
XemyXAepWd5a7J/ui7I64JqJ6LOcwDn2xKOzJtfSH03UgKOTsBmWutnIhG1KrGH7
1EX7agsLbu0jT5xq1wajEKvXb8Fb0/r4nRsx7hdoZMYsm3cd2KesilV/l7N9sAgi
T+C6zAuQ500x8VAZHFz8zXK139D/dAHjJFra9XzZxc/vAsZFbX/y3BiwV90aKks3
57KsQIbzcGkjgKWDoGGxDGxGjVDhyUF0YQhUPy7GyJtEkSGu5clVOypDzUwH3EJu
6RLPeTPVxg39gI8DjeTYvW3FtSuUztRVDCi5+/gdo4B+CcbaPiiaGzybkbGzKamr
IMwBBOoVaQvQRD/quS4U5tOCJQdHN49ecwonsvJwpxoUTrBdTpX37HG7cOR1jOhb
oA4Ug3hmxP7ZAdP3vSgnmdWzX2TPicYdLm5YfgbU+BabpXcW0kKdmFFCd9NgzjTX
Zh4pfVM7pkjfNomsvToWIhwV1oHlK9Y1z90e/INqEUvsWCjglvaa8rRR3KfKaCij
KGpBXEcY/ruTPYL0VsQaVhKDT5F8BKCo6ltediDi7S8=
`pragma protect end_protected
