`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o/RWAAD9ddHr+/+KbJXwYy0AnPcELY0DiXkw/0MdqN0WO8uEyDrVDUi/gRVlrrOf
ZQA7XwEB/kWGFSZsMHx+qrshSjbN47A1NN00uqrlvrz3G9JyJbo1Zx2l+Wvdl6C4
zX0ePGkHUv52ySYuKqAODJVtlDjJ8//lB0wu2UG2Gbw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6432)
USls9JILzWboE/6ED7jgvmxTGtM6qIzgPrac7QIS9+nY+pvJdqqcBr5sgdrEPol/
feOvbAiYmO+NYEXXZiJPf9gJEeW61cJCwLSIZflYvcrl92KI+ER0bLLBhY/rFpDi
k0DyBtg+Vg2sfY92+R4T+5+16bSvwzDmg8uG3M5mg403FfC12Mah6Dwk5tJBhXHe
JRoKqnDfxwG5hE+auqpiMhCXAIbP1VKFnUA4+ZVmDVGHG5pFqLmIPuv+xxPdqU4i
aPt45F51AZpf+nTAfquQc6WwRrfd7qfwO6loHcpq275pWNUCOm+N+HXOHbvRz5VY
+ZhyRvk74bxrqloK49IjxPxEPJZ6XoIUlZm48R025m+igtyBCUhBu4v5ePQ0lkzH
KZ8S79R76Vxq8xQ1f4cra5hk0bi/nnW9Jmc/wmXv+mYaOf3dq+chCxyedcpst3Sh
lCo5fKypQvyHjR0ET/1rRyaaNe2No2yJf8NkFyP3uo1h3STnwBjAHse3tMkOg3oS
L0tzb16E69TbCJSab+hmnc8yRvQI3W48VbE/O1PQnw2lYv0HNIYgxhib90ids86r
UlxYugs3Z3OymJDmXLkbV/te0dohArgM2UbMDJVkssOwQXcT1yyBTOy2DGNYI9Bp
zWmYzCzRI7k4igN0zACByOOIixwA2H5AuvwfNpVFVqS5pByZzkAt5i1njPFygSDG
pdqUDJet+vJeXzwy070idlY5+As2TnvNEaolosQ8A0WbMln0F1Wh897frIbx3x/E
WYGPo3iut2Q9YZ4zRUTpWyYPi1WYIIP7m7FPlpVDleZw7UBm956jvhgPfYSJffll
n84RfTppr4XzdS3TVQKEXoSXD6yZr/8Cgve33ORTyrM3SP6P9ekpi2IfTXvcNDFS
Pi5q9W4qhd+M9OTzkvxTpjyvNUbCojBdjJPgP3vh0aZWPR3SklATYPlHJI4RcDDk
6QUCdUyX2sgWeMJQkycIx5KfbwhQy0+rQUm21DMkISy1rohH9F4zpBRUeaDn3fa/
LGeuVlkaizWtARCLtuUjN8vpCjB6TcMZUpdYvLDWmkZXRs8KsgS9xUR/WYxEZvi9
9OrAqAFw0Ng8P7MPyDhP1jp/kt5yiG075iwvTMEfj/aP6XQTCdGyan8uRw5WzznF
mIZ8wcmNZKdh+zJBgvMQwS9/6+SObrSmhkxms/LJI+EpcBswKiSqhy4rBJxyaesT
cPOC0JtNoEerFwVZWe0In+jgjbKjhHzLui37iNBfM0XduJfcDr33pD0Ag6F2emLV
xGEPQFGuqsKGjphK5YSN0Ams9NOy0SzduFl8c1xb9pfbRIgLbThnpoo5K15cpIsa
WHHFMhS6EFNAulomuwjCOSCX0tx9c+NVyjUUdmy7xwL4rFfmT7MDsQcNeCXA8+B9
GQSlrHWlj+QAAzFwlHISgopojEwe7I/FwW1hqA2aNHrs90Bx9THYXgs8B0nPTfOq
NTQInKZuyNWaP4YOWgzr/lv6huP3IQ5PF03/fpGTkTPzT+YK57ulas+xskeCQBOw
8xigkj3n88XjMRstQU9wLwEjQ3QPK4qUVff2vf/0YhWzAxwv/mFl3+tF00xgUwv5
lfaO6lCQtP7o0jxDKxXHC/kfSlcFh4EWCXL32qpxHWI6klpmlUG5koM72NtUgoRp
KoBbRh7sDCmpqiOhyIpViATKB+5JuIkKKZc6vhRjQwe1y17tUppUaSaBGtR9X2Ph
GSLI/KDuCOw8GuVtiztnv1oa8A4QCRFqtYQ1rBdGQU/vrkybV6c2ngwoEhKfDS3Q
fMTf+BneUmks3Yoz3tzwhko0jppIOqLqr4e9qIbQJRxXkJ8ZM1VXnEWbqLhB+flG
okEb5ZBW+Oo/J0W8tJbQ7nNRkJQVY0DIEPuXxDXuBjZ4R/N2fNcT4iukFeqsFuiT
rnOcL09kLMBlkkF90qJfqwZ4jv7icfzF2/0Jn9s4Vg06jagoMg/lh9IgidiimAAG
HlDqrg3WpKCiW2Y0Shf3Az/Y5S328TrpiGwmPO9xwk7GUWCfRk5liuh9kmClcVJY
oKV0bc1m2SLRvQobLhqs8CNuWy53T6fJuosK3vG7+kHKzPNCmtp4ILOyLEV0nLN7
OvCxeE7mYEiFSwMDlYPLRy/AqsT3pnKnpDFC8pPjVRi3R5Pf+2oGeRzQkxq8Te9i
d7RDtmCmFbcCBvlxeJvooapiplUzku7xstlCWv4TRZhYszaPEyNO9BBo/enJ3C2d
WUQ1cP2nN1rI0xaTrZUs2qX312hf3G03BcXl94z2rgRkdtaIh8fe62lIjBGdAxW2
009iA1Yk/DlN+aI+2VADr/PyILDw10sCVnZi6JJipGDvpD3UzSR3FajQrZBIQztB
5YGa3b7bEMur6OS8I9Tn+cVk0fp9CnYWRBk2k5i555zKRxwGdqnQ6nlGzutzL7aT
Znmcpj4M7bvwu5j4+VR8UNARjGE8Qzd00smeq1O7jGyAkhF2rRTsXQYUrs4+g9/u
YHD69ocn5VVP0IC340gj62seVAoiwHcVcd+BGgoxrVrMv2PFmZBTZ7+nWEP5fq2u
Ni0dmlC7SOuz7T9++vpNvXV54BPJG6sfWSh2BVO3X6wua7aSd5hddSvRjXhUus7+
m2HXmh3/bA8FsRau7xPC5RsJXE1GrrwQ4I9NjgVzrU/fzNtE1rhzilysjax/a9x+
efJ+2GB/x75JKDk6w5Nl45p/Lq2X0j0kxe3aHK04AH9IFHIeRt5sdAsizmx7YzL4
8qGR+Q0FgpLuN2dz30pDDQl1YDe3R+Sd5xonA8bl1B9mU54R3CFhAIkweFCZPL9O
6hD1AxRnP6qbpMC4r7QPEcVpL+wnnzXz2n7hi+4++nQZr81DenYCDGdoENPZxv/b
FyUBx2B5u5ENEIJQ1UGpj6hLWPFJSh+S/WRhCBvEzxEpYLjPnb8fx9DNy6qPjILm
UuBvW70JXDxwNKOcano01F1ynDyGyGyuNJ0ZG9aBJKH8vhxqsQZlWmenP/9NWJyC
CVoinWFBoH4VgvMm93fArPsCBa7gmGeinAsQeOF+nk38Z02oG4z32+CbKvK+l7MG
xWQDIt6KnRy4iGPEA3idbAV8+AeAf3zno4452EiO129PViP+CLp8VgzmUMyDsFOJ
gG+FuPAumY0wJ1DIXwXrAaDkzzH8lRoSNYzh709KPNz3VLnxtqbZKgaTIBL6hvms
ki1pVU181upcJaSqLY/ZKZuFIF2nBvvEKglvqvCEHlD5gvz8LenLwPoVCGYEvZQv
XkutIq3+Don662InrezBLOGZ8IoW/zNWloTbfBlAvf92P35+ZNLk8OdLw55Ohtx3
/ileWw5hjHxaUEuhLxUKlQZDsCwCj/im0fFFQek4xQrGihTc6TtBojJC88K5qQFi
8dPLcUkmTwJcRvev8vcQOSbXA5UmcKlQTp9IDUATKI/4R1y33CDDeiDLSHNBeA5h
Q8KcdxeRRGXE8wIZbARquykosEALXjGT2ujt0d1463Id8r8RAnOfoG9rKA6n///E
1boW1nHuR3CqhCA/i35zePSbPdcEe+DhGKenGDlz+9Xz/neRX9sz/5jMFCGE3ULg
BUcFkqLslW+bJMaysZKjltyTaZPGc/Mmjjf4y9DqRjbzCCMxFj+zeM/r2KyOtE/x
SWGvpZrRA9nHKm0UGaTdOI3gPA2T7ismX7Uddj/wnip4lObDaFF9jzbY5VPlo/uo
/CKT9JkFuZvSxkkuXJsTFn9AAcFgO0ckjoVzgECboKTbAZowQvr+2hlMWU+guC0y
11/XmrmXckDlibM4u4spg3vqBNrQsA06zpZV1RAwge1lrDahkyeC6cscN4h+/TWG
VhRh3in5TPjEPOwkmNnS6Iy18g86WnsUoKu1VTNcJcH02sr1qbrPqnd93kWM0MMY
w43KVw+7c3GigXttRr69s0pppecIN3A3J2ZMaKg8A9y9pqTIgHkdW2I/XuW5kHfE
xg/JcKL1el820LTGczFVaEmX8DxY0pE/4i3VhaHqAk1fL428h2Hy6DoXgmnMSl1b
EY8kSjcTdv0YRE2hrrONPelA0etx6deYgfgy2LfaG764OtuLluX2beGMFktyN0nQ
5D/snPUCxu83zqw//W8P2ny1RhtWbz4r7p+W0YYC6yqyUFgm/ZOHfmaaMW3wob4y
zpcCLMX9TDfNEsSP+gMpxtQOBNYygw3qRZRubG3Lyf4dKRHGMDIokQaDIhRJja3o
rK33TOE8PQKtL0Gy6urwjtZJlmoERp6isc0vRRVi0Kbve/44PdTeDXHLhyFz3KTl
NTqE7YefBvSb3GJH4Ha4/nDD6yFLp738wz2I2ctj97ps2ktQ26/6XGttmPpwO3IQ
pMiR1LYnW3HHNDiaAj4iakzNG+Q+XaLEU4K7RF7RVShQ/xf2Bay7Yy9IB6R4+uEf
XzKLkz28n1l4y/D+NnS7t8acwUTB+6XTcWB/qBkc5NjZVV4DlidWHoCm+XNkOeI1
F3NpkeGI6YRHPaMWPF9Mf/PUgE7SOOomYZLzkx1XqKFhTmoL5ylsafFyihEOoOME
JvRZOIo3chwQo0+1CV3Wn52H+DmtDfPCUK+PlgJwcrZdZ+hjHPoU42Lmy7kiju+T
ZYzZ/3cVUqtqsWFF3qx4Y6xSIwThDFsatX8y7g4D7OTYc7bI7Hp9fCaNxrP82kf7
KZHRN/D+BcVL6q34AFsDQBkdymK7cTaDLLsThJowXwyzjenMuXOiWShzGHZdVmR9
4Ak2+Es4KfLD93DPCOe2mUknkWc98YkXF0Dx//BGQXIUmPcA0uv3Y6iCIfXiD/be
LaShTV8Jiqd8umVH9XkCLg3mcP/e6y1kBztPK5Dt67b8OQiQCS4L6sAOFKwqJ8qG
34ouhhYfZ0L95+TlzSDYfOcpxOvyRrsn7OR7NTiC/ZFZWR+ECpXxutxwMVEMtPPL
YywAlvOq8HsTK7L4wRGM0bCLaYF+0Fqv03wXQfbmpqCQFJrwhj5OMPDUfI/lH9g4
rmZttSihsVbB3nMmuStNDpj+9+sA/yq7Af+aYnELFvMW2tSlJ0lrJ5zbJeBnsCcK
LVtvbt85knNWDmj1cqfFYle82LvOswskJilrXKPNgMkKSiymnyQRR8X4Ajss2xPc
yhsPH/OY8e7vGxa7FNrnVNVGmcfsFExyGGVh+iuIyeFDV4IwcLZKnnM0jNkY8NmW
h/Cx6m/haz3kct8fZfH+lQANkNcAWVkFzOF1l8l2T1YRKQWsLxwGQ8yxCaRqhEUG
wHKvLz7NFK9Q+wrbXtqPjUSQOflzsBh4ApTBnPiFU9pqIFTQjJCj+expWmZNTlW/
KqoEpxsASzBDf8ZTokceSpUH+SHiHHwwCXQRMjj/U3dJJBM1X0ISP2Vw02GXE5aA
aIAOGg3hLfstFIutcpk0Ez60GvM7hnjOiCkjxTL777SxDgaZfp2xCHXhyQS+P/PE
cDF8SSGTZGDk+oO1Zh5tG8+f3W899YeqVd+IvKM/KD966dciboowPME0T9Ud7Qcm
QTjoNzA+DD5K3JZm8fEYDqTkLjPqzSIvPOPMgCgcYHGpNfTU8/2I1MZAdIa9srV8
mLmhaylA7YvahRhR6ujL5YB99MsUXaP3OaF7z7v2ay9He351vF/BWerNThrNu1pH
HT7Xcm1swKcDUXo5iD6JvH6kda6LwRb5rOPGvf3QXUwT80WziSBU5LxtSnJYOw3N
VY+ajHPkkekaJv/UTEciA6JdLv+qYCcNSLwadDcT5iYgzpS1loRbYoDGJOo7vvq4
aoI+XauVmUoBb8YiKZY36kqdQCRMZr4EHRvu1UaN5Tez3mslrt6z7ReClRIIGnwn
VPdF1gtUiiMCmFIqyodHl3kEVL0T9XgvomEwAqx8vjY9pMw9Ijotu7UeDf1sq+Wd
wX8bSDe1qonBdY5o3OWX4SszROfGLiy6/e8/WIzsEfc2acmokAppTRILsZiFwBja
roj35cTMkWsAjdqMaWE6EzTO5ePc6WwcgFg5FiUeK/YD3re4SnziCuFnqP3RrONd
jTdltsGtW+65yUcxmu7jnm+UzAoApkGaoIgN2knGjBtpNBWdYgynCg8pVxNL0d83
EFMwR5pkax3xdsQDVbR3DEbnJYTZBGvOOyNxlFxjsV3YEKUukVCuTMxu3uZP+eFw
m5H+yewUH0/cWxTKmWr6062EE3CoLhcycZurpXOB2H/kbL10uP97oWvEZzZo2qdu
99NQohy7t0TeTlxyWMhwzmWb/YexFybVqk+HE5baC62XBKtEcIDes2guiiRXwToP
beulbDbNFDPQl2qlI2aCNvxoIM6DbN7MogH/IpptiAbT4nrRfohHLX01HLIc4fJW
HUMXjz2zuLghEBTYr50hP99a7Y/wU9vIGq3aCv0MZc09sXy0+p8usqKy5Zp4hHZS
D3m6WfAaS20D2FCKx6R1PgQklWchoqHK0w/0R1BYb+VpI1iq+Sn1MTE2NYB8GQqT
XSRxohtVI2q8SWx41vSPkiP387EozMJeV8Zr3y641dcbtE4XJ01D5OLnsjXbT63f
6M50Mts66qfw+v9NkaBb+dwsOGhR4O+7jBviy0v29Yb7HE/TcuFlXxz5YxCPoBZ6
MBQyopyXYrW9tyBSdRWaxvotWEaNCp+8uJiNUsU0Qi2kw+XBBlMhbw3d5MzRCwI2
mnx+trCnu25d+xCSSswkowu9AzFaysnZMFiVel/fKcJjg23staHGeQ2YAv1s+sAS
ABjVgNHibPvr/xoL9/5jU6vhk6+Oq7xJSzLkc509uNd9u4GPlKKsCpufWOYeyYC9
nynKD4YTrZ1ZvaY1tjIAqzE7+QHm9vCkcmLX5QHIjleIpeh9AXZm9SA2epTHDljP
IzWqXTF4lTtTjiD/O4NZAJz6rsZNGbFb9t4zGjayhJt9+kiJKzJ+roMvs3Jhp0SF
SExYRLhMtWdj1XyLBREUdEY/jDdKV5uF6zA+wR1J+vG2kpjmq/yR6Jnf+cLAOMv4
CIiHN4k8kcFaTDr+j2wK3B4OOpMXFLsCoI/OS10RRehTUIrQ1IG5Z+ZJC3/ptjgR
1MbCJ6BR+YNws1Z/8aH1LvaYxYIU0Lr+qtCmXGjmF3H7Mwif6ad1ZsMhbXJ8YEAw
dPeKPZBp8Vk5JY/VluwMdhdVCxawB89ZjFkEDzVUWPegdWgd+4dSH2zF98JJhq2j
Jt1RgBHjLk0gFcFmRJ9/u1LuGTwokJQYL+Jl90+SZl9WRr3w88QysltoFJ1bSwcC
jsCTnixKXiCfB8OVYJQM8DFkaVTPqv/KANzmz6bm5mIS/zv9WsKOzAScz8LN5JoA
DgdPmmdZBTTXpb4XQ/sZ0JxnRKoAZCv6Busy3jbuCI9kvLarZ7ZH4rb7IX6D/J5k
hGvP8hBtvcBNEbbXLOhrkdBiUegpmTlTmPUFPhXLvaahE7qlUTmib8dLlPhrEkbw
1ShBjtomTwNH0RXR/BSd2p2eBqL2nTX2df4zQJcAiYMk0klGof0y94N5Cr6fRmT0
/HG27do2yreFS2MKSedelFno99MzOteNqyz3IpPkCLc7Fw39xgl6gjlGE8AhN48/
MyxfqWtbK5rsQJMpIwKevpCQktWV66jl7+x9WmDu+W+GBzDqe2QRaWSF6o01yIo5
f1JwNoCt0ruxAq3iSE4jNEMy0javyVKYm6+2pV1tUVc3e2JeGGNQh04qTqt1ITHB
rnzlW1t61Odck0ypLMe+zyQkCHleS7msgb1InXBQ8g4ICKG+lPm+l3kEUQ5GyrPs
k2RSeHlOHUWUPOWK0FNowhFbC+mkUkdd0/5H622vCj6qNY+mIkWCgBtV/shEJ5Vn
OjK3I5+OEDhfWQN7RNmwq/cuMmS7C2B0bnexu2Akibyxrd5/HybA1WOlXIq42Nuz
l1MvrCp6Cwx79gVGbFLtLV92s9HK/SdhtJ3vKJ2Op7OznMkJpDLLnnnN6twvRsvE
ZYypQYXRBWC/p3u4T7KUBU8vU/08fdt4bOPR6lNBcT/5wgkKUi2XTzDE0su3BvFV
WwusOvRPRnCCcwYDnRgCN3uiuFOTG/2EQOM2NUvxsXx+ucIdo6chQMFKpn0CMH3V
PqWTbXxScjo4ajWjO40Sd/vAyDfB3x8Ujv2DkrM4/5z8aW2qB60uk4cLEpoDU/5Z
ye9DhvHkO6q78uKXjvLJQ12G/v7hA3peBFG0r0H5p/eB4TmVIMXyydW7mb8ylfFQ
bGtVAgj2k37S8xJfvnDKF6v5DHlFhH57HuGtvGN6SRsWeRd56slgemXlzK8g3jJ1
WUPojFPKGgabk5c2Tlf7p/3zIT+Ujz7n9hADVgw+xogd8NFL0PPAZI9e+eeFwPwR
nbTMNoASrQb0T7WLRe7qMH4XmkQNz64i/H0Fqu2HpnIrl5uqhxL54lIF5Wm24cMt
HUYnDx3E6ln4NlB8lLcLll567hLXkVnKD5p/WKS+FRRHGE6Fn71wr4h3m8ax0dxU
IaIGbjgzZHGAktXS5K+GuZ8/3zAjmP72c86SEdd26e/juGExlQ7b0/oagidD6ce3
Qjxq7ydTwVXUCq5vxjDLURO6ui3pK6mrjZQP2UfLbKa07dB+6HE7XPmLKifa0Tac
`pragma protect end_protected
