// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
MDZ5YfiuIoOBLUK1Hwv6/R4saE4abMTyGLY02bHVTz+IaPhw446zfCSyO1hp7epyIRAYOXjFCMPZ
BzB4z/35RSzIjRVolnER/HaFwdFOCpXkdW8Awd8TUpeYRFir0e9f328iyFdqItLfhvtuCw+Rs3wR
RzhRoNmdZrH+qYQFRiLqlLw9KJ6n99qR8Ch9ZANTNN8KsNtbIlEXmB5JH58zj6wu4eQxNuAt8tWq
dQO/kWYXLauvF0+jZDgL0KWD1TZfbxCAG4tV4qvqGNWD4Yo01n481IsDaYii4uj50v6wqBUqQbfw
bsWYOFSMJMPfgn1kY/njkbyVVR6FvWvchINguw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12368)
xUfkNxTufH877GMLZBcAPbk/JSxy303fAJK5l2RiCHQZzV7dxWopAi5qTB5REv3LMm4/dZ6h1NZy
yKC1e52wNhUzhg5rFFq8YfxdNBTCR0vTCPuJeOuPJbg7DNUCIUdHFxezxP7crphcwcEP8H4O4lyp
b0tVarqq2kQYpFrWv3sHpfH1Wn6e5LxxrY2izBW59PZ/4FXjYFFr63CFG0+p8hrG6cmtZZByPMPP
PAYtu1Ixtyg6kyfr4RXQvNg9iUQRVJc5GgBAZeaY57r1NZ53fbTgVrC9fryCln4fRrdqdB0kFs7N
MlWdZq9cljE4qay+W7IGzV2xle+A4Hi0zgCvpGXR3IfDRWFxCS/7uIGoTeBe+5inVpQmhmWQFVzy
0SkrXLMOOI5Hr2KmchFrYpRClJK3WvQ5ENckk6HAlQHLL/jHLE28+7rGCM8PHkRNCuKgAV1AH7kF
UW9HY7KLFFie/ylcD2XMpMn1RTDyKHf2BBvVHCYl7XhPbXMdfFJ2sPj6t0ZStzt10P3Fp0SunTJl
XhksxeDjyK3HRUWLxbKyLYRl4CLhk6r8BUY/J6tlbCKiAEPZcTHNFdy8mVqvBBXDBSTG3hM9+KoV
soQqefGONQbPbnLwLTQiJkbqnfLX0XDHbxFMeXPDTrwV7gBCwCIu1svp3r/l19PowxCZOj6sS8fs
3myTiAq4csZd1OhFdhcKpxfbA6k0ZrlbZ7dPq3kfJ+6tCLMfiL/kIW6OgKWwDMJTeCQkWxW1Pp6H
DiH4G+9GkCPKFhl0KfASQsIXQrjFWD9HE18/Mu/WNqZxNOz5tMbOkSVBvKNciOEuWDmcorpy8vGH
xahG555N0raQh8I6JPmjjgDvjFmoppUSSB27Bbwr7B/RwVQQIoB1pNqLnVnwBCp6zrXXjVTkJBk1
4/tL94gxYED12j/vKyIkgGIodcN18oB+HtqNjcHJG1MlTb6fP4UTVhuxEv3+iCqDI1EAAYeJnp68
5GAtbaZXaHZDb/HH/jgfISfR2gtYIjuJPNhyY0w/PZJ3qHKqJHXAqvDkctGqlZURhFsSsZtgZkJV
ZJztArPEGHyQcb1lxN5GXgenOJ7BMzzPynaEMJfWIIIKYeWs8hdB0E7Rck20pV0/m1i91PIuPnUa
cV6rwfBNHPja00lOBs/v68r9fUXNPjcrWvwnCN4nq30kuMhaGHv/3uPLA4GkMwgkNuTgl58xukgq
Mb9cyhMD8Zmo/DhB1HoDoBmoG03mqCPcKKZXpQ4Uccz78PWOK4SqaYmDmOYkGpStR8hKeBfFt1Ct
Yu/0VIqNTJDpobgBdijdlhYrgU/BqLPrEWEWRLP75U+6x3L/hVGKhr6jjyadE2Aojim5uV1D7I3D
NxgYF2Xo1l8p30EiMM9ml4tJTMYtCfZHX6yyjBLqYd4NtFMhodpcEeo3aLhQGI2kKkFataL7ijHS
ZJGSPzA73n5RdH+YcFE8Y+Q9KHx0YWmZA0Zud3gxzCwG6PGhYlMYYhE4k8SW0QFXngRVdN0vjuzI
ACPBlA8VMFrrmzvHd/JmInUWuVfQ7oDa+RVZHZUi9sZCPJdHmdkRKAlIZlYsjTQ/0k1Ab/SR225A
CWJ8DCyJP98+7DYMdCNWDwb8XCzI+VDwHs/hg0B8FTbpyHa6xSBRKXFIbCb3O5BBGoAswkR6GxAL
RMW9hg1B0ffu8yzDlxQaGKmdkZl68nLiZJaMY8hhSZ1ebZ/tdIozsmb/pxal54Vn7G+lnoEKca63
kANnSxyhsNAJV1c2wAdP7gDpZriDRpKyI7wwi5RUYRIYcK+sDJUlRo88bea7T51eT1sk397F1ES+
ba7gNo6GKrSU6MmC+GcUiiFOQhBmW0Y2wuvr01cJsGQ08LAlzeNFqVza6iSWZIsnxj5CKb4mWKrt
5acMbrGE9wqaonc3m4SAFfl6V6JH+6zoKTefT//hxvF8RIknr7BVMK9s12+GjXGSyRKmQPgri09a
VKnybBwcBqGyoGhaonRiOp7BEmLs7Rj1msJFBC9PfvX5sxRavubZKwwd9ceXywz2H07qI2kvCnbB
3vGIjEDXxywyCerng5SLyfQ5QJttKNF23BJIBgqbKcs1xk4qLTAhv1kt63QKgwDE7mRwY0CPHQn9
3Qt23R95OzxyOySZ/PmweKuxreZ0hvJp+4px/VlYubh1oIFi0A4+kmInS6goAvj++ovJEiVut81H
Cd4lpJV6oDSOiyqKGrm4iSw7kdd351llyoHPeYdnUAphF75BW3vSNKiQeeGqu5O5lZDqOZK+NV0S
uEmWxJac6eASQ+jjWAmkcYBnOO4UDRPdS81EE47ewF6gZtwZ8GfGAXyBvegqsbPIp2NqlJIS6rUh
YZir8TFLCzxEqoXKhQRcEbVEgM/u4WTek9jRxIG2l4r38As+XsLdxo0vWDtWS3lXVhD8kCP3HGUu
sS0KAsMCMVHhzg6l1rNZRO2IFMq0FWbE5jegkXfWHbaDGemQy2XO6NssJDtgYNpxlNxZaHpcxG3F
Xr/rNyltyvBZKJiYEC/ApkmpxR1j1/Y7YE8BfRw/wHafHy9Q7mGZEWE1GLOXQip6PAo0DPLynQ4Y
9LwUJrr+lis4H+nTH0WhPAgfDDYHGogzQB9CsSSU04lqOjtJxGyYvC6TJ/4Ixvgc5xvWRroRn1Ke
JXHmNweo1tb654/uj5XelQSRtbDGoZFRtQavigxzGOmjL4Gi7FR88zce1mKzpdGJd0/jPLxMh6Rr
VplaC00XTuBnwkU3752K6SRhvzJx/QGFrA8M6CzAp3w/y1J1BpMbz/GscYjVtBOoPYR7SFO0p7ur
gXYzkOeHpnLJ7zw2zPYUxZKFoBYMJVI4x4iyoSLpEFVNq2JCCGRHIsCbTVGN4CvafpKuaI0ejNa6
ViNlnK2a++3rASWNQWos9VP5EMkKTOBEp1JbcsK7Eph8VuHuG/N0p32Dngs+mnColhvrE5XAhl2n
MNKA27fcHsyFDO8wH3xDOHsYiCePbtM0N3hwkMtVxIGBt/Uspdl5jCXrbbGFrBY09TiZpi/Asipx
aTtlLlvY9dNy+fqMH8gbOedMRRhOs5TR9AF1iM+R9t5XIHv8c9LSHjKYYggNOfYc8UVBG+VXYO6i
R3CGryjuYYP0pdIWqQ8gDwm4OeyG379uuZ1SHl7L9RnZMKITxYaz+yUZVEKb4GQopH2H5aXYPk72
fgPC8oozuTdBpilKHPNhAtIYDj6ujVfxJ2SfplIYbs5hHH54OD+l9MH6EtFiGmTBIZt8zne449pi
fwIDDA3mFvXunxyRZhCKw8b1u5KFZkt6VpMa8ojqY3ryLu5b9WxT25bol3CTcE8wZszP/P/3gHlk
OUBczaMyB7ZPEndbHgBaHwYOS3KI0Mk1pjjJnrl1f2un/Eshvlq6m8PgOsxiuFAt5UA0W14Cu3no
ffucTbUwMZnZvbn19nSAhgBOvDJQ3MjBbl657zz/MFi5WGig2ZwGvlVqrH4CxldM4HxVyN51hWQI
pQoZHTPWWpge6P4cGAUnBvD6hdZZ9Di6Cjym9ygwiXReNYzQG4aF8cYJFoU2rGwCMd44/zsuZ44d
ieSqfg+MQ2Ro6PUo7+pyhBrKepSDEsfnxq4E+8dri6RvuY7yg6h9cZBIJE/LGQxByzybfNSnKh1x
C3YY3D3CUJw4cXAQV3PkHyaQ8iDqFHMs6XcWdSMtQRWr38zsEmjL2YaQeogBPfx4oKdKU134omp6
zqcynIBLYE+0icRU5UWpOOJjtA49tSgEdY3xQkf6GtUtPvXK9SO5UNIpW85uTEbZKGWWEcJlk/me
IjqgGUj8cec45C6vThszxi8ejekPDgfps344UyC4cZvznYdIed+MB19UgCfE0HVRcmEtqs5nDn+Y
2LT3oKBI2AufqLL20Bm5TJfo3fbs2/gUcdwwrH0LxrnNvWC4a8EK5E2MF/NLTODNvW+An2HpE/uU
23gLGLAP6YDCmQFNdOlOH3P98UB0JZjnSK5mfm1oeydqPXwTfuHoctcAioT3i3DyBcnbKe/bruk+
6RxSRpubdWwE8nCljLYshOS4MAxgfQjKDarnW8ch8+0+7YyUPzlEsnQX2+TS39z0WdAME2tAifUw
sWWjv9M9cLeXda/ovXi21RgqeR5n/h+/S72a53tytm8MJOf3DvV+VsLnS3WVq8X8/xG3YjXuEAh4
tC3ngsObWuPo5yDNUGG2SLurG7B8T8mRgzFZVTJ8X9BtiYW83IiQ1vXvcKbk/PVSx9D0i94xTZom
dnS21D7z6msAvWExZ+smEJe13/KXmpRwGxIBlxUJc++RFkDGSBv9PYXjLrVXw+oQzP4oS5WYMjzI
XnR3T5BlqkblfZs+aYRw6Y6tJ8lReFT87hK5bhxECK56lfmTAXBdtuqPB88Bz3Bs6/V5WnDugyX8
nq7WKjdUiMKZVTsli2G1ubYZdMhCcWyHHu34FlfcUG6p0s8rZCNCelNoj0g+SYGLFVFk4c2zmWTP
yO3ttWzFIBYPfNUbYoHL4HM46kEPEvhTnhXos3zUoLQZkhZUuE/ByDN7qEqahou0FYI28kv+1EK6
t5mLe04SthUCGDdGlXQ8lGPdlUCnd8X2nD3VieECU11RSDdLHZF1IvfksyeYRt5ZG1Lib3DTdFpB
UazU+I3S9YuoS48bDDsiWwt0wD/h3mD9H8Lb/I67FpEqIvYZkQum2gCykWcUjAdTHMC2XgO0i2uX
Oi+bv0REZpH7GMzqVAhMbmjMVawD5rDm5y8nJiZHWN3j62RlcC9YaJL15F5uIssZnqTqvgfiI9Rt
vBPhb0kKgP+cDZoIo155jXTkc3jbifejXIbxhcdVB+0O5u+mTN9fnyQa/l0hRzwVAI4nA2UjoiDO
EA+EtDNddWfxmH4yhMil/GpwFg2dc2oLa8vj6+ca/VjAlcEt0bkWXFtwRN220DQWhB6POgJE1jcj
oC079DDpkxJmyCMZDiRf3P/d2HOeurHbFa6yPTkMU1zHc/hqYUhuuv01zbTGq/2fCYg8ewaBB2F0
Umm06TGfG0CB0shChWIoJU/bPNgpyFF894uDRP0aw6xpDYjALP2GTKM1Zwk7PQchwNIT+aAqIDfY
ZSFp/PURIHlxt6lXtbTmFuUKyJye6sJGuLwt4j9Hl82YPw5WoOik3qgNBtR8VTLO/omoWGVpydXw
rraGOW89ISAeypel11uqUq5kK0xTdAWIAWy3gwLNijK3FuXcmYf0n3mvSYeD+nYkYy88O6rpuGJC
5bO+VOfAxwTm51dhidqJvfXGByg6s/x3YfyFSK+bTAcOvUf1YaA5GrpXVHcmeWShGNs8bjHUbgjk
zhNE9kdSnCmXWMinMcWreKAjyFwPg4E4P1eJN1EJXLUAuDUG46hMeRpE96Inhr1kbecNBRmfEKVl
jYl5aq1vYJFrcGAsWy8Xt6qUd46g1lT2j0DHoKM0FwhR0dacBve4GLzlK2ck3VbSDQRnuzjHvlAw
0+9MNo0+QJ9LSxLr0VhMYZMdkHfl9cr2Ib35g5MqTOH8e105sufX1keeJvdLc/WPk/tQdNRa+DrW
UbT0BK769XSOZGiNJT1K7x3Q0s8xqeQRzFUC+1LKIsOdm87inLs/QxdA/Coi/nE72K+7mwrNeoFx
WQTk28ixPbaPZwGkmUQ8h38WDlCJS3MoxYP4qUsZxtu+jcpKUuOrFjDo22BLftvAWzMsx9OE/yxI
6GU/bq7rR7BGjl6Rajre4HAgVQzBJSBGY7jCe397nbdEU6Zy8QCtOIubSKXZl25sIuPVPvg6/stl
WaU+YtEWM4tCw5dzX/gKgUXMmh61GPBGz8CMkt+FUNCfw2pm2B/GxklL5zZEnPdtbdMc4VyH7c+V
C5yHZEtDxSk5Y9FLCujXS5dk0/fsRMlRUVIqMIYcwzYbZaOXfOGdU2kPB47Kx8YdpORTaLkANQig
FDA6b+kMyS+ArStkPHKSC5v5/6d1nEYhPRStjUcKOBHQpr+MNCG7ZD49FjwzzgDzRbrBLd41jLes
1klClnN6f3xy151ddnlAh1j4mm8NxH+u0ex1z44tSWMcsHzPIJ96DGoYcvN9KouTZBs6d6GWTnfw
RcO902nnRTVfjKJA7qtcl1+a72QPnDhOS8ZLfpexo2okfjf4SiEaJkbYahd9Ace+bhTJjLXkEVtK
MfUZRFhE8knU5S34KNWJzdzDZUQ+g4a3GB6vjyWX5Eo7+tBE/LSZnpExEdO+ej5RoXfn4PMzzV6D
GwUuBg/L+F6qOW+QP3NDPjrn3Z1TlKEqSbkIswv3rJu+EaGe6RwSkXTBOvDmGM3C5tUSOv8R+iYz
7BBlNwQan5qsCAznWkYYKJaH1xs3PFFk/u4nesKmhy0uL3s+HrkWe4AGYbjRBu4xMlQ3ANP1fmUb
AjIpY/hWQLvfPPeRQwYU5aE2fRSVFwnwBz5TEp1YKHqyU9fV1oUeUnGP+q71vDq512KhOenzwQC3
SEjmsh2IGJgPdll3U19CY+ru6KF26ltoYH/Lz+fgu7GG5d3bicIJaNgnut2jbX95vmPbcTjqG2xg
4eeQ368l1JduzQimdx97cCRSSGZJnRzg0F/UjgTStXv4wE4VW3skDOnzijTEP3eVUk77uhJ3egQw
D6nzHtIo21BJ4kvyKS01EU2D4ozwV5Z0Golqp7rCOf79CrM3bJAEGBfyvlrG9879KLXmHJoalezI
BvST1s8s76h20adwQ5rHx/5OLNqZDKCesNXB80mbNhYB+pHgwP4w2cKZJUOkIFDi5kmJHNPP5K7E
UIHY0uk379wzjxH+FCKoFk3XMfPys25ycDNvftci+TN2LXHK7N1aJbxR37TtmfHGv46AjgiOou7W
7ks/jXJt02XEkAOl4kSuPX4UPmqo2vHyS7TilU/pC9CQ2CKYTyd4qujIrfTw+2Ahsl14aGuUs+tz
Pnc4C4UWBB6U2ocO7DLj+L9u2ecX5L0CXfW3y3I1Aq/Vm7NHRBxC0iyw1A/BhpzuguXsHck0OvH1
S4ghHk/NN5pVw9Ds4VC3rjFnveW8A6LhT/0GcPpQxzsWsbTtBSVjITi1q8xblvR8O1iSLHpBt5pz
gDaQM3WOjoKvaP8fBWUSvahx3WFZLdW8buYXp0gvkzBIWRSjCz/7vfRMRVTR98984rd0Z1ufUNAP
AcKQUU1p9Oq6nzSnm/BiwtemzfBMOSMo5c3da3yWSHTrYGYaQPLsohHQvCi+0KBVMcU9DLB2+2A7
hfSNvTBT8jw7E5Wf00BTJK3459Aheqhbc4qYG3y1LLufBdL9iRqDrvGycrKOwp5CSae3Lb5T+GU5
8iO7+TtlJ45xo2isIu9n+kYul3f+fIDaBgGw4CjDaCYnmRyyE6fkJXqo723uIWUhEhJhVVl/7Nnt
tnoWglJdKL3NTP+W0SS2BuqY4sQ76ztu7sn1H3EFBt5CtjNWiWfvhDa44zSsn1k3CfA1at5Gw+h5
vSItO+Y4/J76cJJkGYWFxnj4YzTgoXam2Xtx1KdH2/A38RLjR4p0CRsuJ2XrbAHGEz2g1ZRyYuhH
3z3EC/qBPlshNtjAWn2pLYcgPQoABd+Cu1FdQ3E81Q5BsOYPIBsr0CbG0+XDQFKG7BnFj5Ar/nMI
VzI89HajNunG2RGIX9dF7JhHVQRHUJJsHYlF2WX70Cs9bRCEFrw5vmvVXR0rxUKdWb1n6qZy4F8V
HDnkpMAS+eDP2rpSBmYpcb9tKE4G6HZdxhgBXe2vx3szIUu8c2XPAQFyX4hBpw1InPVQ4zYeX9gB
Ceckdh9fQGKx7WoR0YS2rRBVc407uBqyDpEl3g8dyzfuM+rFQ5wJw28FTrPoeNqtvumVVPiiq6Hc
q/tXF1dO4M1BmIoSA87QZ/Dq6M6d8csn2A3vXEm3e/K0EKhxtw9XoDRitajR9+6ajPHKrHt14gFl
5HVtbbaPPsU46F2VpPOHQ0nlOAGKrcsI4lG2CamSWY1oNJnkvUcuTMqf8uZPBXeN2klijPBb4ql+
4G8RxUATwpfIJ0dHKQKZTNn1qkEA24U6d2pruIzQ5VJ8dkVIvadDelwAaVLidMPO8TqlmliKHGqz
WSjhjwfzVD+42UQTTMkUBrmeE4jCkIqoT+NEYDJuvnrOilwSYaWR48WBX3GOz0o5+8powiT9ouNB
JYtUWkrovMjKitjTfItm/HZ6slYPO7D/XRBMklNzBGe9Jpx3g+S1rlTUCCgg/K8DUynCrPoLBJ8d
vn3x1QwY1BToAZLZmRjRPOKx8kjGlCaOsBgeupI9CdrFycGhV+Wn8TMaw9Ca9YcxOXDJd0vXjrl0
7Iul7S8ta/5MhAQGXrLvHifZTW2wB2hg+8jgjSF2umDfikuo+iIa/3ZkJKWlLdsU8+m0oUyl3Rzo
JRT9MUvZ832qTHL9+5nqM/l/WztF38nhsuwPFXnLeSZpi1z84Bt7nak3qjSjthOPu9+lBHnKGYC0
suUPmUn0ZEDZR2y4HKq5NynqGLMH9yHPaU6bxgTyEbVLOwUIhdHcOSveIVabBc/P0ieEaOV7GvW1
QwLQvrdNml3wcmthTBVRv6RCfS0g++eDRziK01Mm94sk8i6ac9BHsKCExxBfE8i62r7i+H1cSXR/
B2XZHGlDSwGABtUJ4RAkygHV9Z8bVI7gFZ92yU8nUM84b5MEe+EOuB/Gj+FuR8KnDMlBpuwKlIpf
sZHPDKFEg9/TpXCgvjpaJnrK4+HaHvbx6lRkrzsnE/y428kAH8phjT+MfekDUIrBxIHEEge+tOT5
ZQeqBm9xYUN0QM36tUrnyKE8m3ngmEPlEFNM0/2QKLWiQhi5A1O8y0nQcWe+R8AN/DF+fCn376ly
m5QqV7wxhie4aaejQph92RCSXrSAvMy1jdwH6rsVgq12E9wmMnOFI5poHbGJvYoF5TdUXI/xi0Xv
ASRPv9UyZHqPoUmg1f2hWLEVxxOGgzKX3gZTEldH5gqiD7jHnx6Jc0rNwLLMgTiSFJW7cw1x5TO/
fDu01qA0vDZg4qhxf1oI8VfE3iDxArQhrcPiH4531BR6Hrj3QdttaMiEIEJdKCx5x8vm/luY4U77
W7KWfJY4Xsn6Wck+T0+yuBKgo3DGghCm/cHeaqhJsYyrn+bWIzRM0iOBrGQ/Otobn0KMrNdWfi9t
JCQf9NlFGnsr5nd+HqzOL/kthn68CpNVAOlDRHtWJKUngBGMsx5Gk0DASdUZlkTlWSzoG8lFwE+2
lrjO4tlIrDfk0kYRviaGj1GGgLNXknjp1mtIkzMUx5Gv2HngBvr4Mjf4WOvAQFWbi2A1Ry7RigaF
5FHhmK7bmcC4/fKq7VkTZLQnpk/4m0ZniKkYx33boVMjfh1RRafNQxK8socax3CMUR2EK+/+lnIh
hYb6n+SPGvvwdjk34du+zD2nr6vZx0aFn9LcIt7Aaw67oJZDCSi8qZxRfJwmnf0pnXbgVXsBSOfJ
gYzoJT/BMAZd5I3TOXC6fdCeUuUw5HPx4APplV5cV9XJHk1ObQIrCPfNtJ075n+Cor7DUl8d/0Jf
Oo2jty1k4KbFoO1ZW7Q/K6s5lAj8CQXYy4W1f+Dk5CDyglebhYYS6/d2cTJFBMV+6MZRNZ54zx8s
WMH2ok43ERwcXUqtrOCwlHtVYGC/+AffDZunGbU2gjJJrd6yWo5rpXIAA/f7gfcDFVVbx67VyL1H
n4yTtyCs8pkWsxiZkkMo2xeVVcMDdASjcdDk3/iDpMl0zXlEUZhL5E4ckSspdY98AHb52iTX/mHn
55W/0wclREZQeyj2cxPkbpgUVSSmi7dsI3uff7Y21hCes5n1BHts+vaXYlHNn2dZt8ndnq9NVm0c
Cj4eCJ0Rek3K/1SI4u4mZOc+5nV5yVXNJTPSJIMhw2hrwszloJvisAdl3HWQOrQErEW4Gk2qRgVA
CPM95yilyVRl4Yer/MLy5TVH1sn5x+/gue+4gAQq90GxL65rJoNbitiuJUgPI9wmo+fqVLHX5MJM
ZkNb3yfPvZc2O2+jHJ0n5+/JoBkjzbpC7ScbOqpZ+FTyiz+btFAXHGpHpbZhE8+ySw/dYFnyySXe
mwbbNmQhFXzd3OfkxMhODUNucBaOspBOxtx52MDU9dXdCcehB/HvwOujVaqOEZDVDUvCpAE0kFrn
zcX6VAuy+7K9K0CilB0z2XXPJpwPLYCt2YzYGoiP2lozp/Fa9paPhLhn/ejz/VYNjXzPSc6TQF2h
Ku9KDGAPN7Y4gaPg+rAVYRUOsxqxNvDFCuZLyYIzl2P+tr+vyz4dLLjZsTm84w/7v91HlBWKs+0w
uQB7lZDk2jVURlSQE/GRtUlYet09OlY7v59kf5B9TGWAoYVuFY3qhVjyhpPU8PMdI3DvLrRRu+Hr
L0VcZlO+qVx0FjuAupu7/C81krt52n/mpMU3q+un3u2y6Zp1bC4QvDSfE9c/WVs+xFsJwghAzjJ9
SbREJOKhQLduaGOp2v4oaEf7ySU/jv48pUSsNqmR9JHKIiYAzfvAU5GT31aVNdA7A2hLGlxYM3vZ
OcRpyxZldZHnlK92/i2KV24nEU7SM0el/kjMKpUk1heRWGoqWP5KjB3aENPW3zzj/aQl1wOFsgTP
QEl4mIC5iS4J8JeMrRV2IIVVtJqNCk8aqMR/HNF/mSFPvX5uDglNDSrMyBPJtzk+ptOdPOxb2Pat
rPHM80jQK4XJdgf1XmWoq0R4Dx2nN91DY88Yvqb2cLwtXTxB7ZorwBt5klGr0onyM15UfQgUuifu
Sem/15NEAKULyyVHN+SC9jk07htpk2oD8kQrWXL5w+R0G9GROxeKm4AaQdRa7BaeabAZtN3ha+Fm
1sXRcs7yJsjzJkbRR34ECT24nZE9IjEF5lDy+69B1KQ8Mm2W5+mqpZS2GkkEh67JsUPeBfQLWc5q
QkZE2x9xD5uxFw/iEifQrSekp6VPsjeR1yuqEMRZ3+IFiweLoE1gAmyl0jvPvGTPWAS83CSVQPEo
pnz9NB9bfgp6pJ6/bXDSc63LBuD3s+aNH7zlc9ZpzUPMBkNYp/wNu56XBCgeyLV24Wp4E9t0z15d
9uwEiY+rHxdvqVIKBNuWJYlJAUmYH4eNnnrpedr4lD9OGzD78kJIF+vJ/n2dVhV6vo4qHXjT136h
ZEltieMeB/3QKtY4rGTWfIV4mlUZbnj4jXDW+K8F5fMoLRqGkqKiWRwGIHdCznRFMJOa56GJgkgz
lRP7wgUL582DofkwF6OjuZwv/Hgqwnxs4LejG4NeXVG1b+uw+wMGECveYk89AWHLrXw3qeMlzUPL
Y8iTciFLnaJTqNudOfQGR25W/bBuum0NdLGkCOoPRINITAqaqKoPygnkuSRIv/1mOymzZxJHT3NH
KORJlKDzS5kdYGo/fcCdWIM5dfTe293YwU6GQJHCLh9hW2kQlVhufTzEpyNKOUefAePFAmU/vvNn
//N8+GWLzwWZ9zC4TnJFNcjc50lYDRgSRi1iQI68pBiu7xp05Ilf5MUFTdNOTDzMdqPSV4mdxp8O
DUZTzbx8COXKhcV6SHa5IwpM7nKjdiJZFPKdAg1asZe9ssjDmij6y/jQjNiOnBZ84ZRnWY0ezZ37
JYXFpcyMMtIugjKKG+c34WOmZxfoP2+3S4rvf/eQgf4UoeIPAawi2zPPvOVJnBGcCYzuhCXC0azS
0cUE+QQ3zCYItADO1n/CrjoxNlcugnFAgKA4rp3pKFo97loXgW8EdVl8lcQ1/atw2VAZ4Jm45Ue3
XPxSy49oslNFTrIbvhFzQj8DYlXyoABKVWCVcaLrEnB8FneT0tL2fBMfYLqZvHIW3lriNnv7U7ZJ
lBfhX9E9D1Z8TXnfCel5HHKm130SFr8ZhhJZjk8DoHbzMkZ7bzwezxk9BA0S4xPnKqUOu6o4R9v6
FffgcNEU8VErRm4VBW6bEcpQhL//zl/LdcIiZSZYFJRktnA7p1pv5t1n931z9CTFLJiB+nGkbRTa
UlklIe2YB3uGXUQ596jEi7oa+sG/+D1qBdtJkTs+o6lB0C1ByZqfN+k3DIKHNczNWtc2usFqyieu
yrCTh157UqjR6DcCoFYnRFe6PzQo9P/qS/lOaFgKMdfUpH2SVYfyNDshb4G/w+YpPtXNFRhDm6a8
mf2I+ipKCZciXN5Xi5Jj21F73y0zXN2YkUy03rAj+0vFYHwG0/tjfLi7smhbK4+hD/FSJZ0gIkPv
PKOYNoOAtHv468lhcKiYhKQthGq8Isj6MWC9FcxCmlHNF/umwjEjBz/W8Eyz4l3JuSFaIhdTQTx+
4cTPb0+pkgt0IrE/SGMpcYDFdykgYA2hX7rMAG7gcHpgeje+Nqd4HLsJP20C4dLMUBh+XKh/YX2I
KTGQ/o9rE7SjUwXlkveXkVRk7WjU0R2X0lN/TH4Wfq+pJQbWP2BZocgI/7I+o7HN3NZcPFpiDc0t
wMK57yz2XmdAhqbyU9nDn1kGsXSGlOcsQdU3JRsJd9LvMz9qUgD0Yuf75lizr/8DhcLvBOpTTTvi
+VGmy45Rf38Kvh9/uqL2vnS1ib1Ke1k+qdX/5OoO0QXNVa2OMhjPcaLygL0vlCkzuVnJMAzQ2/8a
WdQIwRKNcR0qavd2naAcLlx29LuASdZ2CHrtr43DgLSEQ8OSmU3NgVBsp1+Z6mIC07p+KESmpo7Z
f7tM9c2VyvnLcd2a/au8Ff9MYVIvbgjsQb2ARTNqT5wdUklrVNb0as9aZKBYIj55bNSes/MnD91b
Yfj8YOobiDwmcCVuzr3Y3s2hZY6xDKPAIWswHwJYiZh3Rs8/DPK1Sqvoas1zCrXxvhkfAZkCmFq6
XlDA96IqslstCPrz7gM0ydJ27be0mk3PGd355O4jD5BeQUZ00sBTqb+cvBHBuJpn++fr1rs+jvbV
/y91vN2EDDHea1BW641oznZVeQfIZE0DlIgJ1L4eVqDErZfcUILy5d1JacJjQRhQ4m96VyU3a39A
0vqHSKRUMaLfWRjmNaL/Ktfy6JcC972vBCiXjol5FNQfOYQKZq0QfNpPbhE6MKw/tmhnMEBtpvqG
VLxnIaQoEh+hofkrTi7VvEAV+FC+bDG8TUAeqrwZngVJuEXN/2qc4x+yB/QYsKctlE9+5H+QqfW6
L7MliPbsp1RYMawnfk4+YrDqLY/9tJjcoXW4smLS2ooHQ/DOcZVKFe46GCvMX5/WltFfAqHKK7iF
7oK3nypG15wM1/QhuAyExlUzN9bqvlW/RXquUfvLNy+UuIrbM6qNTRnkG2P0qfSNPOfWG+Xy8nKO
k27MOF2QcPDikZBrKVfXc0603UQaUOwMRVwyLvCqFoQyOgu5y4mAejQQEOWfASmmoDSaicdNlCwJ
dv3zcnRC3nQVu9oJApdnCd87Z8kuq9Wtdco/Pp253FCMVxBO8oW0yGfYJHQSxJCve67T0GGc6bIv
HV0iA+bakXck7/LaAirei0PpT3a9I9W4G7vCsZ/fVspHGqg86p+TthSaj7GlWOwOjBTwNoAMqD8l
X1+EoTUvQrT+R8PgIZkd6G54XHJf0gg1AHQDiiQoO1Irlg1Nyhw5AgexPysndohlH//j/JqCd6Kj
Fb/wR1bxfqj8TF9s2PgStfjtrNiUcRQ1aGd3Epc3U0PieZyrhSy2zZsuLDSSmnx6AUff/P8ld1nw
YWhZLXf4plFzSJ6VKYk7OOum82DXwBaRidv0wc97mh7YL/TsPHhS/zcmZaDd0aEelXktsgfSE2WW
TbsB3bc/Dzy+/zomnHU+QGGbMdaKLO1R3xI4dNKDPT0B1dmbeXrYljZWQmRiwhVmAqokm+yGw+D7
q31NI/ibcB7RkyZ0zu+vdt8TbYAJrpvb7u3MeFxjsog3DlMcPwEmdk5+lOOxBYjgZtIc/xP/KZpc
M9Ytg43kPWEIHOriBDRFK4EXYpIPv7kiOmaiPtplVPDRqJEBvo2dizxCc5YK99UDy493A50TnUPh
Mt606gXM2lLhfJC+c1FMGvN1ub/u4GP18TnOxa1jwrs3WBHFLcnKaZNlHveLiyZxexs8bY78O7Yj
i+u1MTzM3AP0UKu0UthH7x9xjFLet1ItnobFn+7Ke2vK1HP7RTwFm0ZiFnJP7C2H5Z8bcTud/Dq5
8d3234hSCt7+rv09MHtkpxd3BdfqiMj8TKJH75VL9E5byCUOLNfhy8jvXfLOSlwsja82+WWZv9Mf
uo74wSyc9S+4MKDXQYUYlRkeS3jq74U8v5yiQ3VkKiiY1J41Ovg/IG8lsyTydRZhkNs2KmeH5wKm
7Jm73v11ANzPOD0qEJmBxNSBcN3H0Q3IBokCVsX20pJn+FLklcn6gNGVmj4AeuNVu/JpdxGplA7d
qzwiig2rYZMjrRsSxDz7yw96J2CNhPLS8hVi6iOov6J/8I7BkFxJlA+xHtI8q58c5/MZroGv9KlB
xcoDk+jx7ejeE9HlAsyHabhx5p+ZHVYNYX2AgTUfLwtYmXUngjW7kFAKE5+0TSfhFOWUBgBRbcRO
sRZyh9xqqVNwFd2W3G1zK6WmzhtD+mDOGZPqmHNzk+NCKYNi1wNnaLLcy97+NTlbLyjiMqpE59hS
EV82mM2peZiibPPPKpO37MDLCXbTCbvTOOe2d6pqMspfij8K8ogHZuhd24hgJT7SBu0bAyHPDJn3
7gfxFxoyp5XiWX4Yr4nxcZhsjF8aVpp0JLoexybPeAkL4OsoqWbhfY/7qx0bJ5XkH8pGNscjjfH0
yePQYE1Hfda+nl7r2DJNvtVAsiwFnW84SP7Hx/jFjwzOsKkJYoCvy3UF3KfTl5KIx1MuhK7jc/h2
9SReoX2Eja3IKzsz8jCGdXhPWQzYb2rYDcOVcWKn0BjTmfioJh5+7uA29l1pRFFxnNNzxeVxdKWT
ZZcZziZqn4iUzZqYoO18cizKdDiA39aCE1jwIkHyGbXYe5agd5Rd4iABbcQLZjOI4MNqZYCX8E+B
wELhsdM8jAAucj8lTAinmIv8+eAiLKqq4pqz5E/PwgG6ShCP3HjV1V8U+ZEOd0BWYw/V/dI042Fi
BR7UIxWvSVD21oJuCIS+VSc0+YjyWHyMERoJ9cfL7vz9sHCXuVSRXqeKU2k2ZSlQ4WexWoXyIoyU
w25NZZlZdQ6gtP7//PfVQIeDBccSknfRX8UN45A30khMZdGhWYUh8/45aOcL36oIpUGHYdsAO1sR
tJ9dEHEmPMQhFDJioT+1H4J0MHPcH9xslnKTRVcTy+98fQ4bpsm7DirXe2dm0dwcIIb6LSKfqlyF
Z42Nm+XqDm6otoNXdrN/FoGmXKnUdgPyPlQnPdjEjMXNd7+LGYIP63mc3GG1KioBDMH2aqJPwvz0
QVufH53CVP0JzNrHUdmbF4VeZgG2w3+Y6+tdYMaVaKj0q+f4CfxlAy/NzDphZXlmeawZfDp2Nu12
e0fcaU2kzAGDVK+YcfS/ZDHqZuGJ8+OhEq2eg3acBW61h48QnoD398lYvlQxKc2cvxrAmBMDZTCX
2i5YR02FvKX2BnO3DMLM1kf4lu+UsEgD1K+13H+cbsOQ9WgYePCspnWz9G0/jfAQZrCg/owjybWb
bQnAc+9yKSnbs/4lS/Okbp24O44OHVB4rYgSVAOt0BFFxdPkEV0GJ1AwkrjoOJZvNQTIXE+u38qY
E+z/MCOk4l39uFtHYZDyetedf2O7DP/9hVRp7UTkvr6NWukaMO8ZxqEHH6hp0NJf5xES2dMqVeCQ
zUSF/42NFvmnCfsnEuCM0g83+8zVFMrBP8MCufuxH/tM9maQTW6aotnEbV+NIOtNH/t8IsrADHFY
qDn+x/qbbqZN8XwH0UrMrDwjrBFti2HmH1E3L366vmTkMVcczmmVANCq4bPt9L8t/yUCoZgkF3B5
htmy76eMRMu9leO8eJ8KEk1+wMxymgdgfiGtrBfua0BuGl9WTvumbqiEbVni+fvokcOaw/HmvfpO
5EQtTU2aGmC3xb8I/ozCPak0eRFLIG6ScyxDzhiTCPtqeoVS8MnG1SNIiroqZkcmwkvBb2toXw34
A0p8H1iP1xC0XVSkvzS61RfcxSSedhJa6ssMpOJ7cMjhZj2EnQ1LrIvi6QyaOXa32TJBhP96lN2G
NHG1hb5uoQxVli7/SvxRfdg5Oom/r3Ak42G7GDjsgh+IR5PypkKqzOOrGdySW+ym21DJCJZnSFO+
tPZiDvE4/631vGwBQIAD7y1enmpTrY733XSMF7HTrAF+bFk3mbGT69qySi7Dza5LKRzmgkS7gNeH
pdovYilL1+u9B2YeOStVeQAKO466biiAT3shbvQ0/ucWmU8DjiNCZmV1Uppl5KQo4A91TyfTRQuo
FWI1MYSRYEJ9zDLiBRDqDkFLboyY8jiaY8dY+IBt08zE9DQ3IH0T1HmUELHpWXaWlRjMRyxpoZKZ
OjjrTaeXrW5c79sqWtbBHSe2u4/nzAXBXMOfnFiYFAk6tRXHjSH0zShkI3NgJ8sKNxdtaaeQoumZ
skEkTihi56kjUb5r86VbFu6jweaAY1AV52VWRfMYccRixHQpSH2d5zPIapFnlO+SzPn8F2uhoWA=
`pragma protect end_protected
