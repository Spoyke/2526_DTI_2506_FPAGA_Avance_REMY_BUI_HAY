// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
eMrN2R2gtW4ym3b0cr2eVWorls+S7UjnRLL5cG9+X/MgrJ70XCA5OQG43Eq4asZ4jEhjISO3ANlw
Z2w37VffYSdQyIEZ2I5mPRGeB/pHI6W0mBCZ6uGstKvfPhryTk5M047E0mFCQJ6Ppph5TxBKFOi2
OY38GitCggpt7P+88yrl/R2olbXFXSCR0u/eVabBzfcLna9T/OKoCK5P0fOEj+Is8l+wUUAMMAI5
LkRExnXq2i4ILU1Aq9y+NLb7Gk/AdK2fNFGZrEvX6K3omzYjcON+Vm+2/BXjKuVbcn80o2p6Scny
Tu+FM8WtQDRP/AlXRzuTgPFUIuHrCsXu+6RIDw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7712)
g3iS/tncTcJKDr4iyATGKc5nqxDxQiUiAA7KEeAAJj6KZa3cqKSvqKaqM4/dC8sRWsb8SaxsneKj
boSW+lZApf9exHnUboJRKQLeumiDg1C27XrJ0xqyYEdip9pmN+lXx8NNwDkvb0P84BPEROSMQiMK
4zhOehU0m6v/Bo6N+sSsgKqhL4Ge4+IFe/E0riPXCFlZFcHT/thK8nvKEbRgRDbv7g6lD4fckBNw
4MtHX+jUs9AEodJ9DDQmjOOfUyXIt/T2YPikTdJqSVR3xS0lz3M51n4nNvAn2DX1PRjT+K2JH60+
bNN8J8Au9a7tO80fi1BeMxcI1CAEpKa9Ut3Fu+wq/djM8zIGXtoc59+WwsEEIbro898myq3vhBgV
Mq8c1qneUYIyiMQd1riqrCMnmze29F7AfP2ZaPoS+T2ChVCMJ3Zy4B297UCAY09d+3N1S5Sk9xZm
ADYHDR6VQCWGHru59QuKWzWj3L5vtdfOksGltISlrR4DU5DgkCZrLyRRZ0Sm5EPihNrRunmQzkzP
rya1zSKGG95+L8g8G8VcONuQJ9QDSVeOfafPRWlUktfxFH+Leo8UtD+5Pb2tY/ldKqCvvr4Po5Po
KXCxzaimP6ccxC1CnYy/f4OKf5kUpOFC8fNcZlVCed67j66sbDKLw0zWgDbYKbdyyZt2ti9CpAUo
VsViBVJgPfmykA4FJjIwyocZ5KhwoSChBF3vjwWzXhFTXv8Y+zw/Qp8ijO9lu0f8fem7QurpYKqy
ryG1TaoomS96j9NV8oDzzbJiY/FOccnSh+TKpNI0TytLB2viNeoNB+oCtUwH/ccUsHirkemhyEmX
etnpNNy4+EfClfvyqA63HiwM/F7En8Oyopte6WBbiPAMsQSjItDGgMvkZQUfAA8l1atrgx6pBfW2
qCkl3tkcQp3zxiWLFsDIr/6IGjPlupgoVESq28clmJkTATngZ9tzSC0f46fBpregbf4duD56PHQJ
JiaQVO8FZk/G+tKYrapwWap+LlWqIRHuYg9zZWYbiDGMvuOniaCn9tHQx6/Pq3ESgfgSQyAMeaBk
WVmp829deFLOseeMi0cW6oD4+OWKkmfEUuQ2WNTiYJgOv4im/TPPAuWclgbQz+9NsY0Cm3M3Iewm
ws1YD/Wxv4TCetEJ8x9y+j9nYVJBTlBVkiwfuTIVPFbVrLfWkehxBeB3cgDPrlBRSZ5BlZOfAbhO
Z/1aeCu8RgN5OuQeCNsQ5/5whOOPibeh8lRejcL/modro2hhTkJAyCroUKGfqDt+EuIwLSopYKan
epJ8EfML4IpOg2d27YAoDtBjIkt9+5J6d+2vuLK5m1bQRVO9l4Ze5PUjIx0WWgoUNTGizWCTAY/2
YBewhSNdoRp33ECb2DdvZueTBaM7IYK0XuXRltTzoE0sJEG90jyKglTBt4ChuUr0rVFih+/AiIXA
3TzguQhso3CGVy56PfPSqsXWc1JruTqTBnYplJc4O+ITnI2S65CFafG9N1iJc1NhCnqTvxcnrADR
1WgPQ2tolE19OVyCvHiJs1ozr4lQZ5S+miX3vJVOVIS2KuC6bUgb7RQYZcNBUSOLRU6Cva9K7BAi
Vj47fh5PW/rFggm6uH6/FE3Xy3/z+unbP/vKV09HST9HMh5hog+UjLlQc9bBivmpdIUkNmC7Uqra
RqvFSvLFAZsSee+ASVSBG1c9XSQWUxONI3VZXj8Pk8C4KA+y+h5/OtVdSoWEGKPj7BWe6D8PdNlo
xJrSQZpxbkp3C5oDYdlkhRzB2NfY3TyFi+v+Q9QY0achS5misi2SIO8XPGeWqMyjENgqwxsQ3X1K
Eg3xygXmf75O9cIMPIEQpPa/QFeTt9pUKAf+yhTnGeCW4RTXLEHOeJ/44HBWhvjbRnXP/xqG0AIp
RRAkgYIOcSA3h0Rvky9F0osf0wYXrJ1e65LEE7qs5uVBxqFTH2FazyVaUf4LhEJfQuWFS/1dlYrM
utPNSMJbi4YNieo1wqgyJVb+v54jQW0Fv/dVsOUz89iPV2RgpDo/DM4Wr2o+PFLT2fB9x/ji3hcK
XbkHRsTDtA8KeWfqR4zj38lEIvMHN4w2wi/HVpyvQLlOjeCyk1goXwoY827i2LyCVQoj5oaZWlzi
9BKNuhERlTTjkiYSmKaBQkLtuh6iKV0DLyZHHkeS6fIa9SFB9+Jo48JGMBJ+bZeuXUbRmbaH5Z57
qa1jR5vDBE/XGrEt0qMEv4roFUszzuhPTKYz3T+g5aV080plBIWVVQ/2aZ67SCqpla1CoDxN9b1l
Fr8UUY5H8bqth00+LgVAHTo/oS0WSeNw+lf9HGIuxKfKvFA7bsmuitNGCvko5DDj7vLN/m2Rl2sS
DoPo+V3nTucNUUC1wTDlUtpi57GXal10QJHzLCAn4BpIB6AV3MteGJpHTL+feVqWvLL2I9OP/YvL
yHgk+W+ttOWzJEGkBYRvlK7b6yMswt3AFhmmI3an7FqmpH0iuG7Ijy7BLJZppSDMJUMOoRB3rh4Z
DlYgER0SxYqC1M/+8K5pNre0XcF5r/HPyngjKXDUobDhrqcSBFlJfilfiv8EN4Nwl+MI9dozqaj0
7Iy4B4WuFDPqrFW2FZ4L8qAU44FYqhWSlCUwn43chOZZ3vO6HWZ+0lC0AtlWXYiYC0BwOGO4iv3w
osHIT/KC0n+lVAkwupdn7nMWZi5FjEoDwhU7TgzDd7jozij6XRZzRgw+APtZD1E+ssWa9WLi95Cu
Nf0HZjez9HgHCFGbmJfbEyixRbC6YCUBN4TR9mrcGLen8F+GlT3KpfF82KD7Zdy7U3uZXdFH4QCQ
/tOGOY8b9oZAN1UL11qeM5uXTLXYesTcTeJxMMHBWj/mWssv2n8RD8EUb0npF83vT2pds5x5v+PC
/EwaffuAFQypG3fQOxOLbGJvzxT2tcMQmRc2zbdvkHFBhVJiwSuYdjB38RUnv7/oCr9w5s6NzcMr
N+S0ClvJanpxYL9Av/CJOn9QtRRHgemWXNIpCkizC3FormpZMiY6dZJWRc8GPg8/yL7sdCtd7Gxy
ahe9b1qmfRmgDUmmAq2WtaX7bZQbZAS02LwkGcKUPGayK6Hyqme+v81qbovRpDFjKBEwFdv7taSI
JI5ji5xNAFfVNJTP+mLLSHYiTI+FxNACAWPdhju+A2dHa2djws6NsLXkR9GfUMvLX/c8vb9a37aF
FFMMeqT87LmozYYp5gjJcOvx+wJJxnyMtxb5NfDtkFrdpAV738+VE8BuDw1QJ4pSzgVdtQIqv73y
P15/topYekctiY4hH10tx3SsznKUDuHA8Md4eoadlkYUR58CVEgdApYBAJ7ijwY3qS16j01lgcNQ
LRlWHpkEIT+niUGCGa6l5zVAvU+d43BER9QjwQWMni7bBGD8j2m2I1wJWkmNCq9RsvXqlNzq096A
hCuOsXUlfrGZ1inwm3O8MIS206MNq44cjsjDTrrmSPG54wff1M4fVZ2ZoBVLFKaxl0EIPu02/Tee
EyfI5thn15wm9APsQY2BcEFRJ/Y9QM6nK3RgFOuuTc8u4KcbUDmeDx8cEUlYlm+IEq7b16Tx8inG
UhyjKGqcoiitCuHNImCa1vbsONI8Vx83IH1InnpoFYr5et1eSa7Kmxz3WpL2yzaC1eH+KBWhNRqU
wqvr/LH2a2iLs1G5Am1f4FdV2xZ6s2FTZNChJCKqbWt43NUfPF3BIilgGEcipmegDYf8lIkiPmHC
zQoUK/uamjn8jrlhqlZ8VJoU0EfeN0gtL3TTfztcOokXqyuij0r1q2EPCHBIAyeqCqfaILxViwJy
J6f04zh1YQgJTrA9xdSxiYeBAqSseQNr7oj4RiFuIm7e0e+aPobhZtdRr8+b6J3V4MWQXjXfcv0Z
MZu8WWpJcTYyDURbbVMjlr7dj/R6/Dct9otF1GzAf4luC9Am1bx0hG0CN2t0u9XxxADyfvxrklQ7
d4g4JoWBAOIxLjQhY7i2DLdhv8gcAwRQ2ikjSjBs2U6GqqhyD4EtG4+ZvWQKFnkkSqgZ3wYYxkjH
klz9tdeCSPJMg9RrUVIX8mln3ks/Zk9prSiWQXfBAmH9B9ZbqX18eDEq5FzAvOUMOlFmMkhVZDyN
BxMzQa8/M6M1yijcOnWbloTnGYf+SGcHDHXnEuVD+HHAxiCv/z+lNB98zaOmwsVcw6gv8POvDFa0
W4IZ7G7FGGEWpQRC9dCLYAL9thywsFEbFf7ObRhKDK+fNLKfTHr9VnieXUbj2Mj5MZXM+nsH01cW
nzcApUYyHdnXjb8VNqcBRu2MVFrbjx7NuxjiV5o5bS5EE4sv9j9hBEkaw7k9qB51wsLH8p4aCCKU
MfHzfv+Gi4eKoM4QNNpW6+GdJUtM/P/KbNNkJrvDvFoJOye6W2XCLq4YSkMg0/RonQMVtEHzavsD
RUmMXTFMiqDQ+Vs9GwnKxie+hLzeyZNT3k6sCHQsGuvcONa9PHxc+CcrjFugSn9Cj3Y5vOlQkyS2
8J6vBgl30h+IG9WM3qQpAotApYj3EJ84oAYIKsnEL2RajPrFh/Mq6v0WlsxKvZdHNNPd5nYmg0mb
2k1eK0igsnvxWx5mQs8pLKCmaUwt9WNNeWOPVb9Um4O74r8+miIKMjHLbdnzMaPDd+wuCiA2dpvW
2Qy9IeKKjokRTkt3bMypiGK6mvqjDUga5vg1H8xxDaaqPvqydYkqBanBZ9ViUe3ZCh+wRiV9Wj0j
9hCBSTvPfD3yLGnjlJ6vbLLNzrF5ZnYVCdxUSCB0LwoMmMv6DdkahnZDu9Cn3cquZPomqVBfxai+
5SwtyxnXclezj1VxciV43cyh1L4f3jiDgRU1fAGIxQttzWn537PL0ycOT7iRJsRcVkB2iCEaLjA6
aQpSfWwVE6nqT+VJw0xhSv9+m6UcpZ2/Bkg17V00gPK8qWbMZsdmhv9aHuDksxweGdQzwYvLc/OT
BU6zE54How/kTscKKXE/YjGqdcSQhdCdZgmWXOMHXGKikUMFOjadJmJ81kJXLPyHpUkBgyjAlTKy
Vuz4UppKlWTM+ar4ZuAyCmZauqNk8vhM8LfOK0wc7OL6s+Uz1wqAuJ77SVBBWlB91bENU4Um1kuc
bO50tfSwp5XZ/VblFTmac6B3Q59+7sMMjpYh4EDND1CC5AtXetSYo+z8TI0vUiTG0Oc6GqleNpgc
kilFYm9DsM9/WXY8R0Fx+V0jBzKkV2Ocass801bn59Z/6K7CuR/RqPqdoKgylaTgP3N7sQAQRYFS
m0G1fHrZrwDlPF8jZ/EUMXc3Pl/woOd4P0NG1bLCaAGoli2LHa6evIAXKFOZx6WCexHxXONCzfzL
BI6GV/Cl9n+Nc7A57JxwhVTkmcDWq2HN/jKcyKgQzjDqofsGypA020mcaYKDS4ht/pJ07YcbquPF
Lno1Zu9Az/g4jRMswNlVBc1cQEFqtcHNogymcWhp+WeanJOqXNQrz0FiHXiT2uRtIMCo9b1TWV5M
UF8HpyRpefg5uNjLgrPUC37zRF5ZFu1fir4FhR/wDby0i5Oz/k3AJK1aRRjmpPBeH6h1ZITC3rYQ
aZqzvSJFgsEC8eyVk6CSEOJxR/lqro/g38iBrqCWfdpvQm7cQ6f2tcm51y/eCHHH4hrK8EdDkgT5
QXwI6HRGm0Czk0XQEeVNABbVJ3nFpg68lzrfJ3RyU6ylq0vdSiMCZwfTnkuVLdZgBHqVCdlCLlI2
A/7DUD+8x7Cz6+QBfSmJXDdFDDwbzfa07WcBWS1NqRRbl30XtWlhWNyaPLtUNV1+WG4tzDdkMvH8
s7oJzBpe/PpXr8l4Bfx6otkXVtw2YDFBbYbumEaZz8iwDsMBnUa6cNh563lU3KqL7pQ5srYfWkMi
hYk9UPm1XyhbJiYiHVSKdOeOVhxiMgwLTnl8sF8S5LuIAumDvibTIXzaKP0QjGj70wde8poqGrEw
BXMtWLu8SINT7yxTtiU2DT4Zrk0M5Im4ihNeBpT8tWYY88Tdue+AXvll2KqrvkPkkw3kWE7pgL8u
6yOZyK1GucIC7qJkoT/NrSMjT21AlCKF4OXZgIb0o5yhpm2z5Pmv2UdLdXOPOK2bsnYC/wg4jhnm
5JwQ7X4uogqYsYXruLG1NpVJWN5Xlpd/HP5vj/cuAGd2A7w7pYLXKQtC/Q92n/azj0kkMi/28FXi
2UEXd6XSEtDu/a/zSjx3K1jX1oIHMYCySR2shw9uZal8oTO9asdC2ON0lNWHbG4TRJYE1dZ3m8bM
I5QApno9eoOW2kSKJ22b0Vn8pYSS4XgpphMfC6rt40bwUeY4S0dX07Yey3/5hLdt7Y5pFuPGl8P6
BYrg/pCkua6pTl2+Jzbee5kTucalnazHseUluMEt+lhDuDEbtUl5HnRwYQ5Ys0ugGYykP9QwkuaJ
YgWEahy+vjt2NJb5iQsKtjmvyJfoeqtDwYBzy7cl6B1Mz3DSQSOBwi31mIShZ9A6T9m/ec6oI9Fo
pph6Y6cvG0y6GYzFDqJDN1o3mF9iPIAhHyX1quaZCVkuBlga1Dt6oWP5+hDcAZldBS/gxJE5ELXu
DQp17A2Ib6GVyHUHge34QD1uhYv34IaY1KBdTDL4ObnP7pvZikuk3CQ1SfGojJhlyDzKeKdWQ+sQ
bUWvP7zEWYhtGwiazKY6R6cyNqLdX0AqqMlOiMwvvwtbJZmTuSg86KHA1alRVf6eQjsIrlpgmYYy
3ub3ax0nppHhLmGFC7FZBJTPuXJpYgoUxtZMBacDfkrcYsEoW81Updlz2Qk7bJZB5UvDvTZ/+3+i
ktCfF9Zq/lrCzoIivVm7BGcNdSTPdjENz56Qx+abdGgSRjTiTZgwSvHuFuG+cbKmOH/+kr1AkBYB
+tgN5VyX09VkpFqkcRE9/cjxRZ7etQb8xERUaIOGtT90dIvOLg3oqCE7PdJVtPUNDGf+90LfqV3R
0ojaEaGORcOxmNceDrkDeuF4+AiNpxRCMZHpGo10OK9L73j5pM3r+/3V3ZJJiuP/7OIHInHS96B5
FWVh37tL5vWiG7AfSXnT4Wur+Pd35x6uQ7imCPNt5YmzFldGEgnD9pvc1mA/h8eQcLYb7r2yub3v
cFAg+rIVBkMIbJHH6flMDC43fdzHrWsRyqBouSqsFmLlv1rKGYqC0X2L80EFOY6l/k1iX2PWZT6d
eTTpmPz0pbjPj6NbsE5U0V4r63WiBsofmAsW1NtfytQPHfipEBGvmM+vnxmj3ByMG5R2EdHazXox
xeg0v/G5aDH/RDypuW3NlY+o2xwhipXPqssTwGL1rGA8vsIknRr9Un82yVzPWoo+I/k787HiyKY9
vCgEKYhtiOvZ0LnaJDItnIV7Rp1anR/uPLuw4mJKlB4DQQbTEoID9qWy3O/GlcL5oeKK+yAIlRxX
tdHAjEKFyODBpYKhhsWDJhklMAbid24UmKSRPAGgN2jMQkWhi6yQSGIzsk2OxAwUHYbQxzxJTMvB
T8JCtkGyAYKyMf+BGOIHZjccWZ63fcZEwZ1KPAAi1ZfR7oKqhszutX4obmJIsAiXwGuiqIlyKyFT
MmUVbWnAdRcSOdmQXwZjvySKYO94CMX6+vMtcEzJ0Maq8zpGmANmOxAJQnaAmCP8hojb0Oam+8tt
9zB6qareRykQFmLpkx+Di6kbintz4yvH3bUtstlNp4VadvXvJadzM8tUR0r2EFGZlelDLz2l9O6+
gK79tOv37PqrRYlYXIZdX0zwIGrXZI2ptSZYXrLMr+bCT9RKw0F0hQI+TftVIrxr7o3cb4+MZ3Zt
u0kBPH0Ec8Gw3VcxqiaUtaYzKKcLAUV9AcIyjEvlhqtROu8fjIshf1mCdFrCYL6cwHQYJTyU2W1I
8QuIt83cjpQ67892pLABc0RWDoEWn0Kt4tvF15nM2CfNTxTay6/ETeLKrLxZbMVvN4qW6iq5+kNi
SY0rKRFQnzoij9Z8GoTuyHu4WqdqMqcEQ/z6741opoFOuJeO5EpOqeCRyIkyxZTLoMNsuQRLFj33
JCws44Z7rRDncJZuxNCXoEUbuJAddssF6aKFGLDOaKYisyD0kwAUorf4bCfXDTqqHU2yalCzHAXx
1RqaB/y6epbi3Y+3EJWmkKxI69Is2f0BPwjEtzr8ZLmIF54zFQRn+JaKZBCGsTeBedoVg++NmDYB
VAyQVsT3sbADOZy3YWN6h01Z/D7No2KnozhmLoKPp5kJV10vMPL4hJl7tp2vnw4BSOOtUzYIjupZ
XeeM0xULozrRlVlkvMM+0g7SGupipOa7skjoNQhHM9FvUc9eE6CrbleJiLVDHLy0Vq/IiMDC33WJ
zyEW8JK1OwILlpnosecWGEGkg9EtYMWtrbcEWJxU7tG4EdpaWLGf9PVRhPYVCSAcptgymDrUSuD/
6hNoP8xgRibeTDKO7bD3R4wQPGAa6ws8lz5v+xx/NoKy2SluxSIyJw2INHBcO3//2JGH1BxTsvci
1lGBFFX+x80ZLUpjl9vBcpcYOcPuBscE08VR2up6PooGS0eO6Fa6wxfJ4Qr05fMSb+Y+CBzs9D5w
Bltml7gp5OJOSWZPeTd2ccXtwORT0OZKzgm5PVvJWrWHvbmttTkrQiB4dzK43hW6TQNgGH3jEGeh
IoFAMVNugz4juEHFtv6K+S/6CAg4wDz6jpBh4Fsp2CRIhYBY7pXbgOSKf98cF5QqJxo6V16XjD+H
95TdJHHcs/4qRTkOSKa6EeIb6dABmY/u2YkVpR4BXj0qHafiWyX+WyiekiHCOeNCEfbGi8ITXMdG
iinL3VjIQP7IEsN7Oi7QycvHTKoW1aOkT9k4dAz0V7YczFON1b5oJ8Zs4TCKgeIk513A/3KAFKz+
woBc+uppwn4Mq33zZtfLlO3XQN4Nr09L4D6b6dMlfX04bNJFqg2Sio4oEH8hfmZbwabOZYYz/+yH
3cHjXLN3cZnHZ8QzFIyYfSKMq9KojOa2vzNIRj8naUZUfCsTiYz6oeaOW7ULtPbFNQsCNz/tgVst
owuJs+BoEW65kSVYAo9T1YJ0o96fh4zEjs93hCg2N5pelplsL3ENEtlSiQdDZLoE9xoZwi74VgMK
d+C+ORIZFwp6XY6itM6yHqtGORGLzgt61zeNo2avBP9d6b80ZsUPJ8l4yCkJd/1VGKkMfGBLq8j9
VDhKmXktCyEU25TyjOSUFhUQEWkEbywobee0CSue0WD+yhCDW/WyPoGR5RX05mYouUfDbwGUuKo+
sL009yz0FXo/5VxiQVf/aaiueo1/ZBkqgHBxVQrLl8JFqP2LE7aPCFCeZcZDNrWEFEKvjg9ca+p9
oUAG+juRcaRbQo08KO6eMP9GXCe2cMee+4ccKSGKBLgK7HCQGE0QQX/qDIwz4WxJMmnxl4/zRIWh
Y/puYpPLEffbn7yIhca18+OgjgQR1JlBh/eq6fY3kQCkE58ETsDqqPGHdELvrYTOUaBzEgl8SPEq
YG86PulWool5y6iQT5A8bz99TpbBqjvOGqfmLhLPXNXiV5P4qxxIKErE68uZyNIQoPF/JIRK9rxL
meK00xYHFQdnO0mk4dfWSKuuRm61qpdjQYjbFy1qVWr1aEc7sm4bYiI1OUf+t4dzKX0W9+R9TW6e
VQOQgYrwaAD/7n7RAaLgOcp4UEMg3JjwDjW9a7r6K9CRdjoKtEADhOx+BSFn3FjAo8fDUjprUJ8D
hHBjqcQJyFGiEuFORiKlKWIS5x6IlR5Z4uTB0ysgHPpdTMWuJHAAnkZZtqKGxsjVWuv/9DwuQWFF
KY4ewDnWRAngZ9cjPqLSGGkfbx/u6CHgW5yiphrnWQTDIGdeXZnS0p4rUrRCYny59s/sGWUpMF38
JqQMpaBsgqvQ4fyE1f7A/R8IbNNz1ljMzWlAROaPgvlHD53Y3Lcv7S2SiPPfPNNS/4sXslX+bbqy
8zKPOAqUAyey0AzUIt1j2pEJWyDgfN7+8mf2Ed+J3TOGSvhQo+varzaClsR+NEZTyMpZlQonFyVI
pfQOHYnzo1JR7X+sW3/p/qwrY3C0eiPVh9swuxE91hjrTuEqp+8JBscCg9LDqQ6aDYrZIEscndmw
bG+BXLXTNES4e+VI9ov/5pYjT9dgk10Xc3I6FDuluKqL+l2NL7/lDNQHYkHeXnuXZwdacRTsBwTb
7RqtOY1A7pGu1DjRsDM6LaPJMpevudkT2nFeJhW3CVCgSIk3ikDmtKosMND0j/7+T75lw84VJjm1
tt7Je7Hu377WiHtyMFEDSw0yOtsr+q2JD9MXkXgWbVlckY7nG+uaOJLkWKDOOTtnzl2yIWgdyJ80
ThjCFtfkXSe4BupPiXKH0P4=
`pragma protect end_protected
