// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Ed+Att2xIQniNHozb65WkVceu4kxoP8J/oisTYpLRS5N/nR1NUKWtNhCtlJC1vp33Anw1W4/wEOH
8AAUOHQDilXO6iIqvP0k/isEPTDYQZW5e2qPIMEzF7uO4lrxoeEhf9P3GRg9TeiGc4XqOws7J6R/
2H4lQOR6p5gUdjz838b5IVxCDTQkY5t8JORvgVH6Ns0isjeStn9JgOI6GzGVkRN735wJ/YhF8AG8
evwDfNIwiYMSE+A285p+UBj/4hxOijY4RuqHQ7LRnytxuJatXrfS+MBrGnYzFMxA7S3ovesfGbCS
OLlVOumMGNFH1/YXNktN9y3IotIT2+PtNNwP+Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14688)
Dt8IjIyq1uRy1w/AV5tcLzmnB1sjqdZVXek1JoZ7M8aG6zc7v+42prsV6cyH9ldFA3F+gQKPZacS
4HU/IqFUezaZRn330TfyzZJxCPcCSTamccAnH8Fudx/HcGh0xnZSY8cbHZE2ibOqoauwenyhzHF4
2J9zniCEAb1QUQFPpCPAeZhxYNTSJFXXOl1wkf75yyZsv24VPLTfWIpvHWl+lk9o3/yAItm3f9uo
1ooQgUE2X6B3YDQyyNwvpV5XbcaydljdaEtatB4WybFJft+c3p4+z7zsV0qXxAM93rN3RVrvcwrd
ONQSUTltPVEb1S/ELT8FFFt2P+EyubpTOHqOie8xo2IPXor3Pa8qt4ADyl4K9ol709jkYzOUuEwz
tl7ysc/CY7EGDZCz8rJ6qr9IRpm3TjN5tQbWfVRiYyBQIbHRQtu8li5ykPq/qViETAm9L2Bk5OZs
blSaLyY4L2+HWF1Rkq7bopFzMpex2iBSQu7Jb+6zZso/BXDGIxHwSfpKY1npUQg6hj066e+ujfqX
VGxCPFfYtXJQm+5qU2vnhhp1hRhn8/3flqHwfXJjbTUmcrYqgrwYAjYDwMXub5InkxktZYgwtvGI
sFc2vnWxE8ep41duVDWH+iDgbocGyw1g16xGJOXTF1JMcF2967pvJknSre9xb1kON/lQjqnu0rjL
F/6xW8+UsFxhSLwuQVWd/6frl+ZSE8rdIK6atys1SBytnDZ7hCm4VF+3gZf6caQyb7h3orXAj6IR
OAnLlaTH/bM77nwdsMzy8IIv4KiEWX/wQ31R5BrHmDcJWaRIBpdpuHqCwLbgkCOwB+XFThex7lLG
yM5LEo53vkcYN5mDZFLLwwkjKyRnqwkJIqTwg9rIqQmK1BA9HqQd43T0qvD2rF3C6d3uLsw14xwA
BCNg1nbsA/VgBFlUQT8jRj3dL6rnRBl6Mn9WPWIEKROocSRUUe/1GbMubdkzGIvi1W8bwQIhLLGf
Dkilba1AfLZNAAIp3GAVlsvCUCffhgwBH7rsYq5k67fhO07eiaZEcHHa/7NF/pxdfAremYor2YDm
GguI40EgSIrYsZ1jQbOBROixt8VPJs5K7KpgAApOzwUvCjagwhKsrBLgfWL69zkskA3GsoGegb2x
H2DGemxFsy3NmOZeTYYBha90qX1WTXB9x3ZWPHa7/49IPiAdaeVLbF0h8J2sqReVlXErrCZ03mgh
WkgKNrDRb4fjpvv5QzWkUC7Qm5pjXtOcMceI/BmVYghvL6ZvYZ1TK5OoHrAlF436pU7LCuEsYuEr
tq9IY73m+QvwnFbe83bxGKXhz9+EuDw7du0fwMovOFLC6sgdQ55lukFEBJEn04tKDX8O1yTl/Npd
0/Erl5in0GsPLOIL/eWQ5T0qs7FsGsZuIay6hcuUZ/emcSoFWmT7n2IojyG1LTkcmAbUc9HKRgqE
6YqU1f9Zw0qceePuzyQMuBC0LjVCbXfKHUeqpSbfNVCDwPlpmtdUDbc+oCS3cARS+ZojLz7yr7Su
ctu4OKkPt8FFU1DiS9N4NnSku0sxpephVgkeCr4xmf/8fKyM84bN8eoZmhhSnorTjkYfHA6T/g1o
3kY4XBsT9fKNKnwco7HblOBFkQj6eYIQsOO5bL2fyyA2K1+41aBucrnFkVcrC8zOTzkgyLEOttzi
Lpw3wQtOmsfwmBcJtPp9bYrdSqsVxlmtma7ZjdS/0b3MZj6JR9SxYU09cjxCdJKkPWDBSRRTVY+i
XXB/oBloqfeNCK2b81pEhIqspOb0wevWxLW3u/NDPBM0VZh/ck5DtuKPQ+GxdGtOM1/YPeibtoWO
8daBOssaHzUVIPeZ9NMBIytp6Kr5b8Q+rrAorG7G+F1Ah8Wwdgey0CR43W63GY8+se4iC/+xXArB
Gj+Y5G04Jncg09MbSdRRHH+1NIkD+Mp3Hg0XI7DcmfNnyPbt+skg5ZiCjhMb5VIkh1LxwLLI343j
N7PpfrpHzKJY6tXeixzg+zMR4OsY4t5s44fUvQpAz/cCD14/If5e0d/tvmGYmaK5IHNQBtICBW/8
DLWAvsO4JVmlS5VbHq7s99WsL6SrIdPs46uv05fcP7MKsXS8QLlo0pbjt2y4xK4lHlnOHbzVGyKD
31vuK3ZnhJb1Pk3mHJDmoy1zZnqVJQrg2bd7+BLk0d2xqdzwarEbxTp8qI0R35XAuBij/rZKD2kR
pEUqi1ZN+Hr0kgHveLNlHnuE+QoF+qA6L2jhw3JY1rTsWvG8aP/lYyMcEJ1jNciFwwHP4WY4oTDg
bWWu5F2N5v49i4pRamoyPjDoLbDijuyWx+FdipGGortuOtdgoZ7qE66255Gg6kONTBylNhjCvWWR
fYG3rMX3GYs4LX8XvAaGMupI41LJwa1O6VpZkYSGk4xZksAUpq7Ixfz3PcjPHoDEIjBdERQNH2YS
qxonDIpE/n1vlvt3wk5fa4Jer/7AUP3qnGdqUYkSy+hAqWpXM5Ndneh9bTEGuQjd5crL0+TO7tkp
BFe49Pi76RsrsKE0HlspKKn5I7VoEeF9xpcFClzV+0FA7/Dv6z8ZWh1MomPZEMiNw/MGLG5sYirE
go5MkvbcVGjc4pe4G9rB6jOcAO+duROiTsLB6v4Mgk6lZepTBsJstriEjDs8qXJMM6euyY2XUl0y
kR+Dut+4sHM7GgJKeEHtph/zn/NbcGGXVET2du18zmo0YYjd8g89D8iAoEbp5p7BOp1hgw6C9OOl
WeSwPu5orn6rVwKpNuix+/iksyPOZo2LQJanH9Oge3xsbATJ/nQ/uGhxUoA6UluIWPxEI9NgUGIh
WbsA1ybBR1g8kWZQfX8mrUpCwmf7JoWCaCsXeIkgO4S6N+wYTEFAczSCWk9zjrLyub1bGIo8IScT
f1wD6RqsE/XaN1mKfHbjCOuRbxWP6fi9hkYQMYyzUjXK+Ywt0a7kcGBJG1Kal5HPDc0dI1LiIk7D
g90lSoyk3uKOpjW85WxvRa4zBquuM+0NRmvN7BZYlNcYx6c58LgAZvmAxXwY429GsZoVHs55D4Bq
8f3G34tQHjAulfit4iSuhl6PRZfMbunWx8udPO/gHOe7Ck3UkggW6mUNbc+M1yGyeI/9Ya0e8nWK
gN4knyXlwVqIXsaFz/WtROdqRHhY5kvvJzKtz0iodx4HVtnH04BLTvi+Y146TaqAm8blFPMVpV4W
+DKy0ZGdaU+TmSMoNnQQCbRi/UGVoeyzuoHpeEdrwkIGAWAGSTjmp4Sv2pZO11rHAziQWU5hZuZ3
opobZq5QguYdi+GfZnu12uKZtzJgCrh7ISHF9w+ZNYPcSxAyMONX0Zn8sHGwi5lvh2FfSb/CsZ86
/yLIZ+maHBchlEzgbT8YtNPchMONhZB04o3+Ymsw4+1/eboeysT7ZlQC+9RAqP0cLzCeRulhiYER
c/yxG8nxuGmQJfmKvqMWO4rqad5+fvBIRp/JV/D3J54YFH3hUaoIQBw+6AhwkY+CPnA2+wKfWboJ
tpdWB2A24I7fWk3xLgtDuFRCvItspBw56vgS7wxMjB6uX1ogmKt+ZmXpgjZNQVi90TTcrOcMeVuO
gV8wuYELURgej5UkN+BXrXlNFQXthSvc/vWXJcwFEexLVK1tp0vhLBp3jE1H88tHN+GbX3euV6dE
AP310/lZqEDhm1h0Ly7FnqqKl6O6RIZR3c5LjgPrNbi4uC1ZVrXAfpiF6VaG7gYjui/z4leoSf0B
yDT1KJFnTMAuKvqv9p55Eb/TzlR9gBO3L14RtvDQ+pwz4/E4nN2TEAqSwQNfVN83TyyF8eWDwlWE
Js4836ROAGAyk/3B45Oic8ii1Nx9OTLJkXF4lOFGwWt3rIzQTAg0ZynMeAqRM353P7xM63TCMPnT
FSEhnMqP1SjTfF49Mf0QVR3vk/FsUp4628UQkhjpVSSiuXm/qXHTc2l4WbDVnG4p7LW3bGmLiVcd
Sh0gCSh33wsDhMRblkAij7Xye1qXiZDJQI3PE6pweFXCxsujt89xnd1NhJApdSSQpNCBD74Diffc
FNhikJvElWFi7ScM/MqYY1jkRyTC5zoP/i5olylhQ0ftKxKGsQmXYwmLmL5CSBQqXq3E40iXBjN6
M5KX0f/2ngcscd2goiQJuLOHzWA9spOzCeGru02SDJ5+FjARjp7SyPI6QzhQctUz5aFhRmKguUqO
+DEl/PpDt9eDxnzdmnu5DkOYrvcimpYXztRbcmGIN9cNdq2bhucjPWluzabBuw0ZN7gmz6ol4cNH
xCaRGw7TXd24E0V7cDp+g8I8ghmNQATcnYqOEL6zZuEjwKCJigLrbfPwRZFSyQa35FGZlYpw0YJR
hK9GNsrhjz+owd3LmQODVoycERCKt+LMF2HTHprOfuh69XCRkJO9b6Wi+mGpmVgqMYUhPPAi2HKo
OVrBVYSbYTDFGosVGCZtBPYVMO+lI8Sam6qXoilxPopvT5og6444m+N6LNVL5KWbtJqFwHG6jkgQ
xVIYa3UThjQBioMtgsvYo3AVZKh3JuWsGFjo9f9uwYGma6bxjMYvzm5kTg8DGltQTzIu3Npjw4kn
AYPD+/KkZ+pHFoSpL0hvXucAwtWpE69krqCLTAL5N6FGpVFnSDuiOkl964ypMaFWh8elNT4h8aqv
u/Hyx1/OOsdtzbbErYZmvygJ1TGslStm52aFJzS0T192IPH3iSQq78Xq4qGurtMx7y7nw8IcYD+c
Nt8nGmt1E7VM19zknCkIsdDs8eKuLsmuhWy9gT9AsRo/gdwCK/9JNCK/nvz1JucxtowovhyBKsy5
holr2E3re4G5C9MroR7Q8EWBDnw5G9I+bp6WqqVDxrbN5e2thrV6a+ObcrBibKSRaBrKEkGlONaB
am3KLzmlaUmyo1bDl9Nsg6PN1DMh6gLz7mtDvO1oElz25FfcdS5UdyrqJxism8xHto3TXX3C1QAT
nThUNI3vDOSiiw/rmbc+PDc6i+EigWXqI76fucJRXIWuSAwgwiMcNwDG7XbV6qCbeheUrnvLW1xV
mH89LTqZtcmwfSHSo62DannKTZEb2DN1bkhC+ucjZ5MV+TBirpfSSDhmAWV+YHAnPqUShH96yM40
V8QqqThmkprctiK2RZHJXO8JF48FB8fT/Cb/rMVID6MX5UyaEwdRuJTDT1fOixIanBccRy6aXCHf
6SH0Kd5k/9/g2wzHUtrJhBr0USWNxutCcnVNViVwg14A6H44vZM9gERPNcW6EIsayo3vni4bAshi
dUsyT7v4egpEStyBj9Q+RQRvT5bLRL2o6dQwDx4uUxXoBkw6ovvMFOkggQxCx1nxlZ9qJ6UgbfX6
6mZulbDFJt8VfHp+a2RQVejxQFiD50LxyvDIijUx4/XtrFvdKiI4ncJ8qAVQnizxu3pbrrQql5NK
oSt+YwDG+EeS3qXSRGM17L0TUZivq5WMk9Bff2AZILA2IF6lhdh5S50HLeA+SWIF26qu+5MXoMu/
o/F1uJ4uY1skc66oS4MteUUrRohwSx9qM2+yLVS5n+Oy0RltzV7pBnFMJGsuz3P4t3tgUL1w1oLA
rIFCautpqPJNGJckJWu9smD6R5eGJcOtRXz3Y49SwrykggA4U2zLQJ9mMZWvq3KuKAA2+XNkFcg8
TzXhhMYm4STYn9/WKx0oQkMmJthM8iIj6CgZRPiL+UqKi46XF4ZKguMRoUaIkjNGHkuw9aoZO/Fa
XgdJ14Rg5jEyiu52RbFKxdizBP/pxYB1+rbgI1MagU8yOBNAKkIC2r5mBIUqCD8aTakJvPxXUBlV
7KVWDUJQcC+OeqgoZ+N95H4k3TXqTijm7c7iN01ja8qPHFsl4ntOUIE4ujuz6slpteUbcEGJWit2
yzU8lh9Le5AdPzAsq+s1i+C0D4NKP41enZ187V1iYs9GI1hp0rEPGVNizA00feXocAtEDJaBzI2I
a3LwZoRGDTx3WOKmIBVrcBwmAQdOYUY3nscheTvfRRTJRsvT3qD3sKBDTOnh57nkZ7t3w6GxjImz
NDZOdHLPnf4nU3rsYVinfnIUfnMCEyrVn8ak/mEreUqAfJY4dlVOdnaF7USDzPSSoyIJEllpFJ5k
lxKmVOcCJJLvELntyd3rDgRuPk09dleBBR3pa05yMdtUYA7ujxGBhWF+equEj+/KxM7JP4MPKBKV
1OxTDdDHLMoufw2RjXS7hdwzvZk3pOrFTKuKlZwhDUebHNZySSUT8RcfIP7yCLa8ytwLYDpWxzuq
TeQf9/wVDFkNV7oMfVeuUxZbtKJ7Nbg1RDa4OzX1nAcIw4iqUEdytqINFA2srXNbaDMvbk3XI8Zk
B2apu2MCvj0XwIgzBcJzJxK2hy7VsmZzRyravydQP/jTzta0N8ntY4KnQ+5gWxuKRdyeiCtOW2RY
TtqwaPbMbviaqrho+6zQnV7F+xUK2utU4Z74UeQNjHQuV+3/JkHZ8Sy8phPKtBbOlGiJCYPqjXkA
H1ZO3AP7TNNxoHKs3zPPoGem0ofKudr3nedVf5S4fbHEdJSHN4EnZ4MSGlhbqeqRFwlPBfmU8iag
DbQBwc210mL+TedAlP5KjnlXTzC2u5BUJxSK7BAujZjvMk7qyyfuw9K76A2p+/af0b6rnHpz6+Rg
WEHhx3TcT9A5ApJdpcw9x31G5+pa/0ggllkkw9mZ4gv6VGZ3eaYQKIIs5W51Pzrm6T4i2CE3DV8s
ki2tkTd4gNasWfuP1myaDCD2b6kIM9N/t02gDWbvmGR2MLaUqR6G5aWcI50hhGDiK88/a4u8jUtj
lfDhcGscson1ebbywk6eRKFJ/y+/Q7zH4TVS2/kRuQ9Sbz1qkmmxUnC+NHZtBpISLmPVQC6xwugJ
BgpQYZb7sJvh4+QYyn1dmoZ78DEQyRLnI2fnq1n2Q2XFHZjx79qZD/oIVLGLCSoMy6ih1g6kaSSc
HKBocyd4M+bve7LxwOa4gS7WV8v1sK36gkfFhlcWuMm9oc/qCWIhjj0UyPjP6JrOAVNZkHupN04Q
+YrecE6Y0QSLrUdUl2TlQ/xygEbMSsOYov7p0MM8hJnuGX736Z0jahdZBe65UPeR+h1Q7PrnJgBO
53ppwVl9fqiZSnxywK5/Cb+mD62tziLrxr84KBgJ4E5ClL0cSQIpUUTbFvMuohc3J6T5xNMhMg0v
8vzRD79YAruSVnmQqfXoAAFNfIUf7u+sp4oeyJLkl9ciBA8q0eTTbsXpNNK2qg+35qlq6jm1o2HP
PMhyhtVk1ufHVASW3X1DhZTA+yjPL0s3hFDw890lYJU1Nb+o/AE2V5ISS0M+AGS6/9F2g1ZjcJgV
BOTXcb8tM/NrtpJ7meAnxAt43+BZAZ7CjPwCm1IrOP4W6mJDLTXebbNocvzME4QVsN8gmCv8IpT+
JXmwgpke44PIT0/R08oL9JxwnRWHOMNx3swdQQN/xjEGWCYYu6NThdDSuUktF88z5Ig1iTLrGY25
hufsB7LnXQ2zIFP7I1XuuQNQx33cqAIIHt+sqriqpVgsdx79sfpgBEWkOptOatipYRmvNfYRXG29
2wFhJQCPdOlJJl5hUfT5dGZjKVBShey5UULBGYYdIaarT0NPToyfKkfYdZ7yZM4rQQq5l1H78cl3
bJyniHL9Kh7cqYoyd92iDWMYXElyN2CMJQdglhtIcSVWW+iFo0sxvuj7ieGR1rkXdGAQvUjx2c4B
G775680lPLwTN3hIkr7pIF1rJK2AqCtVCXAc6tNRGRSLgJ9Y6+1X9BPt7qOmG//+0EPX+5M9il8M
xkn9xpM6UpjmA8PMAzyL3h0eGNA9i8kZZjTQQDs6ZEuZkbRCy8GaCjkUjU+0MzE5zG6c2B5YpJkq
Tz3q3ZqDTH72RZLCJkcEG56dq7hutUSXtKiP3aPX2MAU+UWKhjhMyVBOzLd0WQnbvlqXFe8C1qMP
FjiXyBXcgZeLIbzK6OPWIlVaZlFKuTf4CbkJn35NspjVZ6DZ7pPFfvut0Jukrj10Spj26Q33eJoG
tbE3oohgAK4l7+evYIKNtfPgwuY09HSQeMHvpE2RaHQMIh1fZM0i/EYig+N84RGdG/wMgbo3bAi7
dWXOaQ+kKGsRJdLTjD4XPQeP2DfeLUvteFnezlQOKVzWdPAiFYC7fD1bxo9N7WQP7LqaFgc5xo6f
DUOSn+QVw5bs1ieVacU3bilicBVD/sT03RgfeT6ftJZtku0GbOM+YLxit6vlHPBetqXtmkf2gL/G
Nde4Z8zGcHqPR7fdEuaHBhyaP+qHJGG2m70QffNpSMsoG3rtBC7HDYK3O6CqRa3Ln/8rnsyvfjix
CRrTPceMYT/Am4U0fA7SjS929VquMYx0G4+oFt7Ut3zjwRVjlrrw42fXSXAQcpNYaWlgf93Ji7oN
Wg0wcyrQHlFmQtrKgQNSPrLqxesgEkT6aaJgq+SAJEfPIGgJ2pDWf1PIGjOO8rPOQpoIdOpvV/dz
k7ldZGcA9GXcZbCXmmmR4laIE2qHS9HF7l70wOPOWdims+E7Z7F9bpBe29X2TRqnxoDck8Oze9Sr
y0X46twkc9q4ouSnw2OxJcFXf24NggI+qb/JDr4BJopuK6hSDJkZMAPiR+r/eYwhT4n1X7/y+EVu
WxwOrv8tdfUnbG4qV1a1M9pGqemeOHOqHUp7Xq36Cwaw+CWVP5honPM58TOHlJe9oOUYdRSPnCYP
b7z8OjKY/TNukDU3CW0QELv0NIiYsE6rhJKOVYAMyEye4+ich3q/XKfYLWqY75iu+XO0MkzYZaHH
ZrV6HjaRG4YPmkeAPiyZndhxl3xyhfz5AVij+UsJ4UDVrt1IJZGdAx5gFAkAqIWmcafcrFId9jOw
65xttQfe3wd6jgt4UyjuKoMGkJeWhLI7jsWDQiGkUSC1bdeSG2iIfE02jApTikMhJWDTO0NPo79d
pRvCM3AN0D2Dn+f+VytfOvst3Pugl0Ou+Te+RePYDs6VgpWk4Dtt57xOQ5xNMKtpKAwKlURcTcW1
F1hDIBWM4U+Ch6VFYm044BZ3W6iKuaL7bB9w180RwShZkKoDdtfyHDfff3tTvO09yldJyprCT2gQ
0Nkh/V6uI3nWdrOVMlgeGxylDEGXg/jcVdihu13oYxPFvYk2Pm8DRwlvkxclK5RTQa+F51zq9m2Z
+k0vEPzhq+2GYl57mPx8fwI4VqV1S+2+pFei30rdb0+w9Uy5ZP2TpTrGnO0SztsKbhcW8NbeT3GI
Cdcuu5UAJBcBSwncOhOMkthfqBehx/l1H5efETQSvSbHkgdJt8rohMVqTKCogOmEYSRKLVbbBIUA
CdRSDRBsQH296l/lUBl7gYpIDjk342LCOf0K1tRd/tjQA5mmrNYp4dsecKgrCF8SC824Y1CK6Cte
WokEK8VluJp5OeZMNPAqssWvLmbWMTZcvqNw8v4uGgiyHP60BKPpJT4ORO7HrFVJGv5Ze7pB19If
q1JT5tMSh42c97lUYzDrQR7zEvg+VjCnVMHqNln8yp2BK24ZkqrnI0gCiuxttEK/POESIXJRwB/7
ugbanvIIN8r23l37p2dMdNomzODVolNicZb/OMbDGksYQtSmy4hQkLCMXlq9tEAQhTb45SPDmh44
0VBPsmO9Lw1Jq2p0Ans82+4p5IgWPX2kii/lKato6kwQcBmJJloohOSAmSNysLj2nfxLeJyofPtp
K2oYovaCy36EaDx+ZokiX969M9myE4mHquuHwq7kdyzu9xI66obwXvtvtLe9gshrUHk9btV/Im8N
2NdZwUIxxHy08t4WNWyCwjq2nTXI9RoSWenAWAlfGc7Wp2rP39Cfa9zWCHP3E7mCzrhnq+59ufYf
yI20X/3iJDfv2jckbW6VMBzXsi7meO4HWD+2G282lwDQserlhu79fqs+XgqhAZqtI67CYTSscAIM
23O4SFAR1rY7Y6hagCJjkVgtLcJ3LM19kE8PiHHW4ahGPwexrPEWLpz9Oi+jNZMvQVvegphst922
K9HV2iEcuOrBs10n726kWyTmfgd9wOx+C2liBvemIcMUzPLuZkKFK2uIa/OjiM7wkBrWF//aiIys
jSj6/4arpDbjS/ZQqf4XVQaFkbUckOcvBTqBadxQWfF/MW3RMnAxuy6CiyljFI5lgyBBK/BrthV6
mjVOclHidrNetFoX3x6bEb3RWeQ56vNyYkyj1yFKt23ZscsVIgscNu+wcP4HOxQ685WBhSiHy8/Y
juZ1mLxqbgucglA78zyf50gUHZvzP/pw6I1w+w6WH7apd3b5utb0Je8/bGvfYGTt+8TUCarEM9rj
E1RxnH8IrobZaDwmZt2c6Da0vBscChVRe3AdfDQ+OzHw1a5Iu8K2yqhJX5V3SndQgQCM9ZPuelon
ApHhxLZKAben1Guhg0rb3Fb+qYTkSOmnfBFeWGuJlQXuWfxaerleoiN8BCEbTASrbl9fIic8JKxz
lCgY9W9x6fxKWqGYgrT2ZaM9TZ/6BoyXVjJbLRZx7XD6eiZLGvIUdpfzZfTcexNapWFkNxSdb+4Z
EpbnulSyrhDf9XCjep9zdmjB4jb1WW8IkRWMp/fj/5hTJ/aagx37Oig236oui2Zb/1impwt3knzI
dGAxuhWQKrQbQYWDk8Nv+VvgqCRiNXiMRUjuagZ2C4f8fem9528eXKZBHu7ddKuKE50rlHJeUdsz
iwixpDMRRq+PzPbaxH3n5Bddv2HhIGOsu8V+8jdqiA7lpo3iIWkjWJ7cN9woZOBsLnb/YCByQ8xu
SklH1ND/9X3j9V0V1g72cQu7WJVNkeVn5pEBxvwXXoIdL0crEN4uFqfzyRe05fS5dgVTya0mZL96
8UL7Ic2AhcLvJMUQ/O/7mi2eqpWN3B/maC/rdYr9ucnQ0QahoOGRnbVX4eJra7ckn89xvk7ug26d
CTLM0sEJqoVaXKRwLyBjt7fYHM8tVzw3hOrA91JkVfAAWC1hK6Xn9IZx6bjonpZXre8PHN4CByKB
R6vdn+bzYY5fn34c3qWeln3+bi0MCxuX00nlWCC1pEUgf0UZ3n+BiqMRGWXueW77ylZU08J+ReIs
VheiQ0nr6DB2Wfsf5NugSdHjhGrQTn1/zmfucKb0imp8YaAaiibEhcxCS1jHplPTuDgri6guWi1/
HqDOmlpn3a6WM856kmipbyZu19pxZzfCEeTsXJew1ndaoCzorUWBaCxkauV39tpu/N9g5bSE9mB7
b9Q4/1GlzBS2nX+Sb7ovhC04FjSAwvTD+tlh4x/LwlDFYLPYm2mYC4gJnXZbXJaGwBqiO9jQlXVq
0WF6sfF1IyaLroyGjkN5dNODBSbuykLCTeqt0KnSIbxjnytxZV8dcd5QdvGeNaoIWit4nVr1IBWB
oF5XhTBRVwhoyA8JOs6I6lIIDfiYP2cWiowYGiiTellvb2dFtVXB67SFfqRruXEWTVx6AOBg392O
7OPPYtYXxNK68eOR+3y4iTv7syNskL4qbr3SKMLbysYGFnolGtq+ZhpDdSahdgh0NQySG9PcWHQl
DQuzaE9B7zivG/1jKvlt74NELUF2eBZeEeTAJYLWB/O60oRFZQSRvAIiPXjXvDayTSeUNSNIms3Y
FHb4VtYNFA5ol2Bf+e4Anu2Am+X6OG4yPRSpcmMNorxturN0MuFaxTjSuFdHfZEhiVMbr0h3yD45
KcyXi0ioBJ3T/pvf1BbwANIKGwv8D7Mk/DPbe7VDpCwJs6kH49gol3da3sb4HiXeOTag/6lbihgP
Ou4L5dRrM7qFCvpiui2sluC6p9DwUT8vj+uXCmtO6GCq6cDYPNsstBxSSm4fw0u2XQv1ZLv+nwF7
o+4qlFIDUkEzUNTNvDF0Cm6VtcwXyQmz2F6q3BJS9IFpelKPSO54lDFjNqCp+7yrLEUF0/8L1hZU
W+xLrminbRH9+xNAQ07B9Pa8MExIhQuaCNG1REoXgDU6nmGp6+RHFo04J12Yk2x9kZZjDJ9SjFDC
f3D98GPiHLJRxZ03EevFa9kuy9b60tb9cCgSqB7dRlwThCznsqPmTReuVEBTjbeDihgpmZpJzkdu
YFFVMxPBxNKIFLgWWUTp2CAfdherPxEPlYhf7ZV/UCn2UprA2WwyEfo+0DTc+vuRPQq4VDeYUZNV
DZhlX1ZmmRnrviZw04lgjRPf8zSlYVGMWbOCX9Lt4yD7zT0s4k8Al9wD17LhwuR38lNTDNiZQnrp
LsmUFga7eIAEg+s2eZAnAYMLMhRR1vorbb5Lgw6qN9ocZI+sgStemUj9TPxrgG+VKGAp1Xb4hEYc
tTIicgp8J7bfobhy3f6isOFR1d1+v2qL6ivGx4eoewYSugMns+lRvnF8PJLk7AuUxJrU+BAbV+7H
ePU80v7PEUkmmAv7uBe+ne8bFwbTehP4+jgPxITMg4XdPyq4qDEpbn5wPGoznRMPtTZ+Yc47f4y8
imm1Mmqw9lhneoEXOc8tzkvmzsrXrcpOdICZrqCZgncrOoV2iAmwDhAAdpHR1xVukvHnbuLHOPfn
YQLO5o9hTQ6PcgOuH1Nk2m3tRrB4zcHAL63UsHsfSm8Jrhn2EOOiZJlPZaPLzFANFL+ecd0HL/jV
Lkw3khsfn0vGEv6zmkSM9MqSuWH2ZvO2FMqqfP7AT1xf3CwfwCmF45SSgDXBA1kUzNOKhrxL9b00
EI/2KxObFxb+4VFH+uzOcir+6f42XBimgp0a3P2t7YLIlzRe/W0W99JwAdjMnJLP1FMl16EtA8D4
wdqUKPReXRSv4/WuyrK3d+O5uT7JzzRGejk2FILdshrL1bJx9nsFKN9KGVxKXIcv0lMBWJPYmR1z
3DtLekHH8LF3K+CjdD37qoc8ul73ePyDRe0AYdw78+rC4QQ9e3Bc0If3W4qDTHWaWpzELEW3UA0l
g4YJtJVpFaCod8vk+w6kidrFd0k7TYmGbGqgTyh3v3nwORzOnsK0UwdGQG85xm0K7ypVYCZNUFF1
LzIFlQ7LGhWTJTcD4IzqO0JKTi73cQNzcS+yZyu16iXHGAcXGU2OcQlDOKeJsCve6rFYj0qgazMm
LNG/L7ozZmuRpuVfSz05Z+TOK33R3pFNO25fTAL8BK6jWSOsYGanVMgTjtftj+k4JVr0cWTaIOTU
geJornfqN8RsHlw8Ic8kD3q1fiQi4l3OdPvfhUJPOe/v5SqKFgHunpuXzedGuFjx4gPH/ox7o95k
tTDEx0/8OuVzXKyAQF5Y1gzn0GZsKiIkzXz7o93CkGORXELie7/N7SHXlRweON5b62a7zQM9MBtv
bmNQW9AdShMtg9iq/EiQ9PYT4gw0vyCCeHfJPOu9D5WOUJsTfb5bR142XW4IT8VHLpbX1t/cmrgx
B0GjrR5xjz0J801fxKeGmp5ovIqFoSe9+RpnKLEYm7AmwSSBwnLnT1TS0UV8zzoiQhL2q1/h2Vw/
nNsKCmuW6MXxRVNx+/PJ7ApPWka3Wq8WU8nLMy4ZfjqAiBZVeloYotxJziIMigJKETKfKK0hKcWS
Y59GZAuyRjbmGZ9uKw2wGePV/yS12NHBseV3E0b77zhVoM8y4YKXgCroFZ+obzNbbyS2hLeFTt3O
1Tdre6pHtrRMWMuYFYKzEwdOsTTkpJAXDDHicBfN2V50S49Edn6wh7tjb9NxOh4WE+GsZ2zeyDhL
hsye+Wwu6yjg/7ECRyhOK3mcnTrmSB1/ERsoXj6ThEKLjrsmxGNlLN4l7VjR08bAwvdfN/Vps6Js
BXczr81yc5iThz0EQD6Y9067YPm6W6BL5HKaIDCDgyAYGoLvwnuBFqYeA/NLtsS10W5OfZoTH60J
fbZUr6Y2w3i2ATOyQ9nvH/ugqKJCkZhCEl26qoAUM709eAS5ITBaihNG4KDil++kuSP97M+O3aA7
/mhunS0WF6krKzDs7XiitFfo0TU5m9WgteVpmB/zd7Aks9ANz0ngpTco5gWhgF/uT3wc3g9YrLfU
03odRKR8uMuPezJwjArMvJ/XgN35dIhQlGA0M82daU6rOIrbfIC+2VlMt2JhQ3+VFV/FN3WDdgBK
meX8m3h9l9L1EdBUKaLG1OhOifj7P3MHcAMtL9gbgxQoDUbB8PV9/Y/ZzBRT0ICKEtaKKBTmjsJk
+MJ8e3GKyjoAtPaKhl14YnGoezlsCX1OdB60vmHmVEWR013Fbv/CC0TX9h//RaAOuksNgjYGuZ19
mkYGHrNdveGeusx3dZdal2NpkbfMpzYlY0PXN17ORikOSGTUQHi58lx2eFv82DoRQXSys/ewGIOu
ROlCXy/dsj8ntcHw1pAM27s6XKNSoCDzSszDLDSr5oTNTm6mHPRN0KhHznIXBQSqpkXaDhoxBP5p
yEoeuyATjgo+MFDR17L4AViRpDJS9XV486Yn/5Ur/lwrqZ7D77y5pevXMUKmahPc9IgBDs9YMegd
WMagV/BXHqMYiIKTYAZCNUJT+c8X0v30EqMnM70y3UqssYwXkW2Tub0dm0agf/jXJxe2gR4Pj8EX
dH/s7AkfDIg5rkICYDK6jULNDXE7JixK2L7dtwnvMZIAcx6YjNdRvD2Iy5ku8pTw5kem/ab5GDUG
+KdspipZ84emZOYsnAjayZvtw942/84yhNaJ+lEFMhGEoJ6mAZmU1Vw2tSOiJZEVm3S/pqjt/wy0
NWqWpH6WXJ76OmxNSXkSQ5dVASVclG3t01QYefp8tJH4pKBiH2qj6SpWjtXobeCUp1xnWYhw0rN/
vkpJ6iNrtFR1nrcvxjWeMfSvb6JiqFyodgiyBXkShyBm+7tV4SR0H7u9OocM3bv7EKzajDievblw
0C5tKBjg0w7TQpQUdL91y68/MDknGo/oWGiOZ9cqVnhxx0yXIycB1x8PcLKpdv1Mh+3UP42KS8ny
qateu/2/MM3RlZzRzuydT51agvjD5kfHcw2tW83lIbPHXKjtCWJUKx1KC1ipk4/PechB17DUds1t
D/+GR38U4OOUWlL16q3kyhf4UJi8qHSzSx1FKPXbrUYK7sLZzd7gXHE2SUY2Kfm4LRtYOToWt8uI
x02/+GTHtZdgjoEG9uk5E285FMmYLZ8mYl1MErEDZAunmOz46r4rXjrVfhjciuH6Y+doN19HmdLr
0dBl2gYzG9c+Ai9/sM7OjbIY+Ux3f1Uyd5zXB8DFWXnLhXFd5KI54PSbCKirCLr3wcyMUZd8hJRf
UO34HmUOZe4zIEuCZywC4mCoZsQhV64HMPL6fUj7klqPiKZ92XWz3S0NfcicMWXbICeqU7MrKmgh
E9LCQY3gc4ActgwUrllAfj4fVZdwuVkD8EdXnZWIcWyBKWthxjzjg0hgsrQD73BYyhPhiyKWeEBs
V+kMzxv7eJk5g4heVguWb6/ytRldmS4YF/6QkcmiVlXsvu/gbM7WOFLLQKpESi8LRD0PO10fJbDZ
/bwUPHW839b5HN+bZNc3ssVrX4NBd+ou38OA7bHUy216nI442eiyGVUMZaRk3REnQ2dHGAV7pZvP
bYVoS+z4igkQrxaEKEpfO4jDG70zgb9ifWNmJjLQAcOLDAVUk1gE5jOUUerNskKZmQm1p26E625s
aePZKDJbtbkCfLqliwORYBrQ4bhypgexKQLGfr6Lx1f/TZRwPht5YPLq7mDXhtcN0ULfuezyUg3z
WWAKmnWdwYAQMErnolhhNIEBmby7eArygn+O24h3eoXiCwIUU/l0CSseh8BJ5isCscZd7ZsFg6hA
6HjR13RatcfrzJDZbe/kypczq8pRQhXic0aQwD6DkGPr7wH6tqEVkrCole7cqG1J4g2oVSjqJjwa
5WxfCav5Mlieup4nOWBdioi3W8isk2iA1uDU4hlM35PwlwpjpKM3BdoGKM5oFRcbYWrwfMjR6ZiL
fDtJZnqeWOwkj+z2J5cOAfyWJ/ILo3UgIm2r3zYiV2XRo+ATGef7a5NQbVqkP3gvFWfAK0MFaXlo
udYDJDy7LpYpyLgRsLsmJl1Ayi/FkWW0MBKSkrU4kCam7ae0TfzuVxipf3+9uxhZ+OdRvZPmBEWA
FXbZxZ5TaUnyuXeUIQbTf8waXcVstHjDY7//qDIfjYOSm5MSdxGNgfXrjegFQkgYirub+XHgCw68
Jqub1EG9B6N5HqZd1CZ0oGbjTt0PdPwyQgrxrOxd4cjaHXdOltb59h897737dgHRB1MGlQdQdaG4
/GXWO6lnXLGBgC3iO39AKAPgDOdeU3NI6kBw/PzZMujT+moVY8R0Di9vy2Xrema9Qeix8G2Wkwjy
nmrm44tkgHr0WcsFTjq5yq+JMSPCRbvq4Anz4wJBIm6VPhQgV7NcLhpykkmzfylrVxA2A+JLxlr/
qYZJwyxH9pRRsfJK31jLxJglXBiqc5zpoiQouCsogr7FOY/W6RY1O7NOTDEHplyFuWq5I3wqi3i9
2xGeX4g9fv13gfdzSCOqPZgVtJfka+VVOZZ3Oao1GFkc1ivUxZrqubNuGh+s3jPICdaZ9Sf/5wQu
6ZTBMNEZo2Q8YqrsRQlMmJ+QlrAPjzDrOC03DpsjNryidrgNjdtiFwbjAx2SV8ZdIsUiocADqOJm
WQFsEBO0EzlVy/jmm50xJ/c57vDcVLE4+FzeEvZ9levybPUz8LPz4kgsdDVtEdEFdwIR7aIz3Pv2
KxOeJ2+2m+015c322JFnVUOsAmH7Yz76MXKwcXmGcaWrt48b3D9GuT2n/7SP61cYzxC+X/VZxwPG
n1qukoNkngbZJrcWUYu55lZrrNktTOOyzjwTOm4OF4KaPt4Q87HuwYc5EFrsAeGX+bqjLVz3O9Ph
uOQOm/ZUFaqCAwc4X7vi/EQuzgrqHXQ88ZcaG/xYngqRBsyDYsLadoRFMIKByRj+wUkkVcr0VfzG
YnnvvYaKHBuf/xrueIWUABeZFCiyPBdRbAHfHqrM91rogHnC3AlIh00XnHnvisLv39NGZsTX7q4D
YmvlQ3WaTYsWM4y//8W97tDonvQuaCCiVcZ2B3sfOgQhSr5kTNuee8JEtFzaSoSdv5R/wF5KETz+
iEUAOJvGPVEKsmW5iIpdVpZ8eK9s6lxUdNqDQOA8rBwXCN9tTd65CjT0wnrp4I3SxixuBUyNB5zL
n5zhhmqfcU/ZyfAGYd78sXNfT2ggasKVAEbAx/bsvUIYIWW4Cin6qNfyBEXALz2HRtP3eYZw5+Dk
znJlWefPs2rZaJrsZGmVmNVzpFcVUL9LSYMj7jFaiNPUm4aBo3nT5zXTJiU8ZdEbUNdzIcG2VYzE
ak1VMUP93yV83TU6plIwt4BL+UJ4MlZam5dLmDm5vUhnSbxdjQU1s5ZwBDExo1xkPKgQp2BoYEKU
qhjNKNPYhJ6eowtrFI1MuGxYcqz1t8G/kA3l+Q4sJ/fGco3F9YH2fVlav9LlcivI/Rosc3+IB6Kx
pPyuVPIeY3BXx9IA9Fve7Twe5jmLlgzQFmrcB7WTW0q+osspWRL6lv7DnOUM71CScJt31bpm7TnW
mHDBEkQTPv/eEyt018C3avrfILndBl+8TmuTyTP0hpHGFfRceVI5iBMvLlqepa6aldY6/yt2Gzg5
y4FiB7KI9fKgVM1B4xlptw1vDuFXAWVWS8Z4n0aS9OyXfO+GbDHFsCXrv3E34Y3UGKoISuswlMHo
Uif42UD+LuWuiv0onmqJO0W/FB8TbjNdEFEENqMhePFoRObkqNJl+tq2HSR37FF0IkvuV5tmmc2b
TAEmHERoVU9f+I+a8fRkfRTQfd0Q6H6hxqRDbq4ICozanLNDDRD/R72vaIyjzV+jd/kvgKpTSSLM
38PDspqgxlj+BOQ30t72E6mnsqoM16dh5r8Wyd+9unumJSxvaEjZPXB2nAqrVj+95h0aB6S0W17L
Fe6fPtUJqkMuwopXrNEhLL6tvKQC9nQnrb6J4YD7Gh/ocdVJpNlQd5NiG806hIir1tQShfUgsk4z
nSPvGfppbZK0qnCQ/rNwCKrDEPrm1SmPo5tpxQ6pl3Ze7BGDnUytoecmZVIG5OYmTHxkr3cEKYDI
xxNTMNsh7/sxO1Jw7JdvLon0nGaGhGYICZGl+iLIAmCVfpXUBPvImXrghrMtlui7nmiNsGRm5TSp
6AOIgt1ll+8HrmySfUvdCA42hj8xKVo0aVg0bkRQ1TyrJ5wYVmyMAxe7037ebhOfKH54nk2ZorAu
jeKyL09kfejDpDP05quX8Cpg5xsK08nAlu2XXx82TzNLCLAIaQtcdLF25XoBePjvfW+ZWDYXSqwl
WGnLTR+hG9p6luftEqrKYMc4+40qbxeoPTzU1Qtz4dlBnumVdpgvkWqjzha7bbMoDdl4WmBXbZvk
tLtOO5qphJzOADf1UmTfA3qdXLWKzmdtCZiiSDnY3CvRiCJHQ2uZIObOZYfS0qgtAs+UoUfbXNCX
G3+DCxn85hXjwqQPy3r5SORUYX9nAMJ4uNVNvI/ZSjsh/akKBP+ynW+9cNXJHjLbIXHHUWGegIIm
9pIBCKro6aUXMjdGCvUbCh5Bet1Gn9h+bBX1ei/bKvRM+RlJyXIFq9oaY8Y3Ctn5RikH9Lu1OosU
M3rPZOXzaQ4DFTXp69Joz7/fDPXYXJyrW6ctdjZmte496i/tCvsf+rV057pVGTyoyX0mqdJ/d+Mb
Nf9Jg6LJrFn+xOzXrcns4fMnbkMNOeCzEjmdSkTXFJAJ/CbnohGkuBribAz3aeLkVJX5TbrBGZBS
FzELmC9oC3u0mTucM020DLEmdgrj6wEWSfQu24ZjBJ6oAm5/NJBxcnX2qOz+R/SsSFFBM4BwUR8v
BCMVNA88w5UH8b8NeiZGiq2O3AQLhXEgXEMapDfQbc3zQyIBhho7Nq6A2pll4qBNdJt6c8K2rbH/
+IBen9k/ZQskpKzXc7g/EDDUHu14fhI0dsq/hKUFJd+RZB0giLfXVbwH0WFdgPBmG+ckRbkyX35w
r0HQTrl9Ve0adGeYEXrYh4aiar/phgex8QN692XkRgkaawJqBHM/W1VRYSe/ZFJNNwf9y9xIvxbs
F36+BobfqMTbZnCI6GWuW++9YWgWHUINWvBRLolfHmG/cKwMkeAP3Y0Oj/FNvfr3l9tsvK/XIgpG
g/aAwuKS8CqVC2dK7cpknznp1LJNgHeYl53TK64ZF3Jc8nD3hV2rbW8KvT/qtg4Nx6JoqVznsOAZ
mhASVXGV7Hc3ScJ6/07xNcNXDDMMR7ffZI0TvlK01hIqAn3sNPFpdXAvlLZxZ5mzuPUjlnECNzJu
EgmHOpMkkln9ufdDQy2i8sT53zTFrjAI4Yzp2VBB3zgSkMIjR4b93DkzGPXSm9/yfDBw6W9uaYB6
68Fd1LVXlFoxs51YEUHcp9P4/tiKjQDI9W8bCH77QTqRK4+w6d50DufBfLOiiXKamrVnbxiy0NR4
K97noceb0iZzHcBUJ0FKIvgUKATx70JC61xvqBrM+9VFQFOgRaD6ide8AF7FCo2tz9n6ie7IWi/s
UREeqdPCQ+Hinm3dTrwrdGR1RxFlGNaE70P1VG2r3kbF+wSeu721GnCxc6/8yU9QDxQEFcjRZLNc
aGZc/qHiHh82usMYeP+bzNqLBvy67u9L1BqqfRWssGAK4BxSbGP9FnKgX+baGAutIQpT3t16Ihdx
xOo2nOfHrtYBhBpOHWfXkfp/4IQSvU1D2AV9Bk3vp0dfcE+R1gMC
`pragma protect end_protected
