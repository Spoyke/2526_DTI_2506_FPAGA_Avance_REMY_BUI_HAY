`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oU54G8y+6vk/5sd6quOyOxtYI9nwOceLHOwzsnKy/wnFA357/Lu/L9aGRYCmnAI+
xuUihy5orGUBg5X9GCILrQHVoOi+SObfLjKNtoxR27gRPMJbZg2QE/3p7CFuXEaJ
oIK3SFzj0qlIZzVgvpVOVwlzoVj5XdPLqXlM5NNUiW8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 64944)
69NRGQMUWBwgZ6Gj/EC0eF0KUpexpmo07VOR4/9ZHbFb8VMd84Ow8Z+iTSsKwKLd
orbCu68mQYNh7utckrUj662n5ptmLhNWi17sHUbqwb108uddXXt42u0XDPgJlAES
qeCNDciKuQjgvXxztF0znh7WoIgrp6HIi03Th0xCGHyoXARa9+WQTjCM/G4mkbeo
PftXsPcuykBuNgJakdxv6WbNHdJgfRjgGRpI8+ZTrUb6vB4vJvnut4/+zKZd1NB8
IlWEZlPxsGKWBktGyHnTf73nqaiyScFPaVxRmSHcIfJSS5sgv6L80fh/XyiZ1GPs
9YNPOZaxZV3sqksv5xpuwOu0KXM0jw9j+2THkRUBv7EwGBOH6mV45ntQcUh9dcSU
3IuXnMFHyM/+Wpit0Mj0Bm2iPjoAiUK0Ku5qNuyu13NQGPL3qEm7Fj3UcA89Ml60
ynLW2csuS3Mo1TYMHJSsUW6Qd0dHTypYMzJ/9qbOlD0ViX2UTxxljW13VqtaRJHy
09n0dx8/BnZ/y7BCjxPqkaLoiPECqwd15CEptfLWVkxp1TMy+xMznTG4PuXjp+Fr
yi619/9QktP6FYzfI5HS8XwHqo+Wawxj2nnbKDvP/Cwy4Vf+qtUQSIoeNqxIWU9X
vbmHotvhxEbW9c6GOr0gjQK9F7RXr/JLKEnWSZ6PqgvmA+Ah21Ecy8d81YiGON9s
HlpeYQu4MrO9vc0pxhrl511sFK3HGjKQcFBDmoJV2qJvi1dZrrbrgoOOQ1n1rj/S
sn/BjLn5r4G79Z5DW7jkknRQaqUfIw8ubpdAhVnHtSKNZRZmOM+oWTRMDASh43Qd
V49faKlRFaur0n5Kauv25T/IVLFDfo07t3doXCLRBRZ9zd626laOPCsoRsyA3ZdD
FoS1XXPldTY7/RZazLtZEwHHgmf01OC7EHcpX3pYFpfWs4Mayjbpw8HelWY3Jk+7
wnvD+93q9T5MJiJIQF3g5FdJFea/VEletPpmIOUl/hTgQfbdW+XIAdx8PauuylRV
X1GcBMhGBqhpdUOUFl/MCRfS2HzUTFDGw16AC9T96mdB09oJjTQdKXqY3IttebH+
+4n+zmGsSn2Rce2Ijzqm2wUUv8ggM0oUrxdEyKrMJDPZHVHwKdLllYbMKsl6Ox+y
PK4qeTLcmFUVvK7YfmMMc/2v0ntXTd8uQSzyzw36UaLoMlYCUK+g9MelpGkidzM/
D+J+VjkpbHVzt7BvlQu9iLryWYs0/OOSctqobJGcfsIxswHuMMxFwcRZJ1i0lgjk
wSr8jC5LgltH9QcbqKuqsKFF2grgldbchy7831c6CoumhLVtFQDrYUKjRb2sW0wR
Qdv7FmWn625jipzN1da9T2ec6AVtMIR2ENRiBgAhuXXTCWXNfbLPAFUB0DRjDRws
EWosafwp58dcLDirvOmiy+kOeWGtsEWsktNKIgF9Ca9e+z94DMwOmEClg3yigf3k
0gFemtgJ/6K5k2AaemLhlhZbK4vqKcpwSd+iiFsSPEl9HpDawBOHXF24OthMuYbk
07/jxx3K6K8VKvr7RWvVRS78CNsO5OXCEI4qm1RctRnJbm8JllSxQH2CdjPMRi3c
Fa67X7LnqKWR4jn0ukDIJQPwtrpKoJRqErhrnHCxbBgmRqleY3T5F2FFvQm82PaL
tL157g6Eh9eRBnJzekLG2cgQSSVEGvmpdgM5ScEJoXxX29Gjb6UGT489NujO/YAf
NVKbplf4FQzdD2BGPnezLyMyhT73SRrexYkLCfOGQtmOQ+LFGMapqZ1940ziqZ95
EEQeBTxSwXJbXflR2cjOs3YMRfrvu4+ndXLCmcktHkePtmvcBMU+XDO25SKQiU1I
2knmY0GwMPldvwohvdyYUKoa41fUkQyQ2aFTwx/+BtjljBnxiiv7iOK5EccbYKbd
lc6gkE/5C3KS3cvstl3yhDvIT8Vvus5leKtkuOPNm5kudwPNf5ntz6tuvJfjHeuS
blyq59hcqHhr+vLIPjMSqqR2ljrpcxEGVW4Ep3McrHlY6csCbltbl1B4qN7gc0DK
0/DBGs9GGsDmYRYZYcn+ubqem8csBWOdAPBGbThRZy1oJyZWXCCINLRqD9lb40el
TxPJS7Y9eRJhP2/HUwKqtfEXvsL0oKIJcx1Y5wkeZ0mPEBd4+4tQDtpyto1Z2B6z
S8E5717CDFXybCHULuuH/QArr6KKANFMGLR/Gu2ilFOEgLg3BzGFjFIQ56mwHaGq
U0+Zb/1ZA9+Z+JG6JAdDXLF75z3fm3Mr9a99tc/xAlzYlq6OxK1saxPPvdletaM+
bpt81trLD9ROkAO+NMel8DRbbI4yrUl5H+MNWEfqWKRERWJCH8LH/pPqsJypQUSs
qio5FZ0LmcnmZN7TPlkIzX9IbHo74t+Z591smyyKpv76aaLZMQaIo7Ykwnf6KBFz
/sEVayaclyTXdqv/pDhH2RKwUz60Nsa7rmJ6kngKtIsAUnEvEN3e7NPjrb+EIZqd
zdzr4bHxcyELHLiMGiiLp2O8c68jb7WOjeeuN8Hj+oNsuVZ3dYlPVCfVLHqXlLcM
1YxBmlYbgThPdGP2BvmYyoy2AefrCQUdpvmX/URsLSfBIrLKZ17rNSy+qakkPv4o
Az4eBbHEACFB1lSmZNrmXaLcdzmaoKdwz/ms6Sh1BPOrN0lfON8LLvw+uJYQE2z+
ylFH/agvKJVDHvoE8M4Yko0fdfSLMO90OY31DmuSBzhm2064QA9tSShAoFJUFzPK
8HXNFCNycimQA0kh0e5FzFzccv2s3AERuKrdGyVs2wcEua5isgfnmdBef0B5zMXh
dts4xGvujdUp95UrHbCVFs18kxOlJKuXX8mvicIv68MErUQRll0wGGQ0SajIxyLd
U9dG8Ap6NfKAcHd1jrw+f44C8eVtIkAmcFajaLdGJudksir0KDPiW94TxkFyeQLa
369h3G0hcw+0FCW6UoQjgKtMt23w2dVcj+pZCxyQ0YhJScMue+91dpcS2VNEK5GE
6/tIvGnmsI3ucFNMHTOxex+gxuASo3+gZ1/LTWo/ioIbj+l7YlO861yqFNXD3SPC
tsOHwDrdLH0XaUUxCvr44pP/4oVu0t6b6g+rNh1CWcZnFf+DxO50S1UNRBVHhgxS
3Ts+YrmmQ+P2MH81xn2IvUqip4UXFWfaqshD0qZGSnlRvBK9XwbvF1qFDEh2jDVh
kJkSarvv4Rw3ddssnpqqqI+iH2o6AikQbtkQppmfdZy6JiuoKfUy6ZR8417v9UbW
psx3OczHSEZ9skBmzF30v7d76TWsXCwIULL/lVPxUdPwcEZ7oBQ6Cj/EOLdebcBT
sRRj1mNDEbz7AHuLh8d537/tRYw3SWAs0ONI7RZWEJS9WWQAyjmS6slADTJobn3R
vlvu8lwZRmin5/1FyXEwGV6Su/0irwMJayzdpYLA7zsFSwM8g2QJ/ZNaJhu5uIVJ
SVWwwqK+XWW7gLESLOBYOzWs1FqTtvOeVcpolRfk7qs0Z/xrGZ6Lx1/N3+6syMTa
ngUNC87l5rns+T8Ai21QiZoEY/yFvMg/84h+bXY04QuCKvKBF2lzBKW/zCxh4NrH
Kwdmv9MHkEI5KCJxKbsFThmZdnZII8Y2HOkymqr+LVlJVA8uKoqExWoDUU51bioH
ht4iZzxze11FRODAB+Bf8cLFRfBO6OmSkAyxU0M3U0czTSPX4xp8TOK94CYK/Ax3
JX3MhlLBgqDvL9LfSmsaINXHw+ySIBNKkx23rPT69fet/0+L0o/aPoK1Z3OYzbve
fTgyzAAAyd3kt4lrQRQXCxUtT2AhrabWmUJFJ2+h5C2NOXTMIDJfpKWzHJDTDxVF
+XQuXsAn9Ve95E4qTrj58IOzmogBs8pWKD4m9rhnjlt5T3yP1qVjp/w7lPvcTFof
E3Z8dIg+N0s4idqce7ITcZt1MjARb2D9FdAw9Wyc8T3indodJE2cv9rOjqNQcUxR
j/7Z4DzLV5gZ7QMbMrenDYUeh9sEtwuV4Xa+P7/fyZaOAKbnl80KVncCYQmKwrci
Zzuai1lvekrl0kniNwPXAuTrekJz28m4+V4AOSctjxWGx1jXhGKCCjyKCJKEhoby
NmGcz2vQEAkTX6K5rbA7wPs+7T1VsGPD4gcdzshKihYIvJAfDbP4s7L0D0P04A6J
dlPkVQDe6FFuyPWJ2/24ZDZaZjPnOcifa41Skzncxo3bPbLdvRdIPeRls9rhYs7P
3xgoTc713N469WLrIXhVch36Tu0KZfmvaOAJ3zW6hgg9o7hNoIneqTgEHqY+QNRL
1vZ8PoGijkq89sWTCue8ahzVq8cZNgEqHREvIUWqjtlSZUDEYcUklw511b7fFb7j
Ca/amp5xmaWjXDlM62pP9Op8OC+Oafleyw8Gay2B3wbObcEMRUnFh/jJeuFJ2pQ0
bgjoJK9m0IR0jyGIqbILnpIjfhGJ6kL67oeoA9FAFQVhMJM5ya/hSmyptL2KMe7Y
Y7g61Hwon2hoQafd3/GhKQ3j1jm3dP+e7HoA4PRJ6C8npotybpruj7WsbQMnKcCD
LjMOgOKubRI2upR8folQa3fLWwMGtGL+ZaLTutene1W8T3uVCXdO0p3W8Vpl/2IA
bQOODEkzg+EFfiCxc9fMwAbQFBdQnB56td9Dk7PS0KRDEtRnX5GoPsRiFbRK68h4
dsSgz/RzzOVDNR5qAH+KEQcht5917ImaBwERU0g9IfgoLmmQNDNugEz9FzQLFsln
r9TAsx5qxZSPwH4TSAMfudSQd32lBOKuYXqrzeuuaD0CpY+9+pr8M9QqjcWlKwwQ
D7FIYVe8EWMrmDCou0YdNBCuZzBZxdGzT/vWpDA/OomVXEhWqX4BMu+dYhWJyIGA
RbU3EQozrw7HZD91ALhz2c5AtP9UZE7abuBBGYV8Kv1C2t47yyCiyjYNrzPtR6pc
VrcuX5xVroPL96GojVWDwRaEXMnQtn96AIOS4IUTP4qzil91Dv/yziSrpKcDCyL4
ddi4JZYBu2x30U7XotHM0bf6ASqyn0KjLKfO6eFE0CYJbX0Xjrnf/gGEgoGvaZQL
iCLJ9OV7YUD4nvJQ93MpzbE5I7wtUgEe9OEE06x2Jp5d2fgXT+0AhVcFS6w2hehJ
MF9i/E6c4WVtN8sso+Xtt1OP794NNh4z1D2UgQcj3ORjYjdag6RLDlDrAnePSgUv
vOcaiDBmSrF9e8F5m90HOlZnybioiHbeLm8Uy+ULhkpnIY/ULRTNfR1KY2DokgnL
yDaM/Qi8p6mrPhkgFq1f4aQh1e7X6NQlIM6s3lF6vRY5U/3oBWNyZsYwA/sN8Xia
zOviT9LVKjCCeDqwnHWISDf44UzQNKM2nzxMr+fFxRkqyKqmh268J/bbaF7I42s6
xPAA547LWXFycl+dFiouZovgHgwymg5KD3F0juUZ5SZaznKgjY7xhhT4lip/Tp2E
gGs7LEwoBBk3diPHcCa7BF7ZN3m6OQYAd98Tc7ejKaD/IAaOyrh5YwfKKrywoHKW
XUkO/97adC/c4NHN53zvB8ZwA1yGPYy45qpCkJPqZbL5KNFN7cBZ3qDx0lt9wDlV
3mZxUzS8ge3XDyalHTbxIQz9taqUF5iATjIl7AnDitN8SmLfJnoGrviR49uiGDJ8
H9CNld2WPBuPXRv/kc7F3fjz90w4z7OsuScffdwMgEm40j1nLMSulFpPOqvtV0Vn
6GCL/kHVa8pIq8NaVuLxFUG3/4oI4MXLAP2SnWdrvxQrrjE2QMlxJm4m0Oa8Kfws
e9mWMzxFF1txqyQKlcKW2Z/NUY2hr0gXypxZqLiZiu2WbQL6sJJvzh6r77pFCvdy
+foq1n1XdtPdgJIZujkYVao2rOBI6KBFn0ZwMkJNFof09LwsXhyOuO46z7Owbb+l
LbQJv0ZpONAYrQ317j5UDX23ppyYcXX57RtjPthwrIR8KZhARBZJ4zH6qnS++Cwq
vr5AVWNjkIafp0gKvgi4M6XM4htVH6IUN6+BtOZa0309EnClfGln3Q6UEcI5wvO+
sohVOPb/nwcwS6MlBEYjndaY9PTdraYTgHKcvH1QOU27Kn7U9mmUlTdlEu66JGHk
8gssPwqAbXJpN+Rn3tzdtZE6PpieKg+hALqQTXqbsxZvw4YhgLqxlY6DPEEfEjk0
uxc9tNaGp9nKU1bTlzRw99inU3NPrLbsFooPH7yAqsU5j5FSKU/lsKinNc397LVb
FShkskB2bWpIuAk/zJQXUeLPgVrOAdS74rIyUp08kwYpk0Cm2I8gRVv/pqNl1Xof
HYeXteQR753zH6/ACaMnBWaS6VXJoKxl9h6FxzS28ymTnhtha+JZnOaOtZNjlm4O
/WGCXOH8EaVVXVHOCzVQfTDAElV+GFVz7rXjK5/7O3Rwe07EVMUPWWgieG3eQ+47
D+wupdZH3NLFnpvCqzJn96OYeEv92DNr3Iij0mnbcb8yVDwjIZR4CkarMqtBzGOi
VYUe8gYtOVX391n5sYkuxEgE636/WB9DG0D6BEFkgy634HJrIEZqVuBf3gM2QRXM
ZUEi1l2/fZsr3hoKQCAdt1QMwW2xLJq6NCTnZgHsmqYuuqs5CpD0TqJg5HCEBa+u
UUgV5zQI8e3WAil0MsWupXf3jM4PtwbBawZLPBXHEesr9Ma4vlp0cHiLCoCRO4mf
QFMcbeKY/Zg3hKRajEK6uN1qdhOezWgaU0lKJjRoGJ2OWL7qlEKZDCMJmEfD+pxz
/FsLwrFcTPZW6M5Kc3EN9LKnfQ9LrIepNe7spXjR9ENmsHTb4/o92cIwnFZNt8e/
NDm4pBzae54u6b2+lZgISdcLpX9imXHPFV1rp9nZ7BWrIYBO4cYdz9QHnNrYVGwB
WuC+vi1j5TKkGxxzt4K0yN4HA/8SWaDLNFj0wTNQ5xrtyyAOCwOaBVVo/i/b+RCt
qk921fpSNaLFeXNwj/Il8f2Yv3VQ5wygA1MetnZJQFiNrVHUJd/3qvECCNJbiYsB
GFoBjUJWiPGq1Qf+zn8CUfQFzZvsxVMYqZtoCNgjKAbNELKFqwrBsQku8zArzrNz
VcomcWDvNLLMxKok5k146RSkWsAPgAu4HlUsQ6kFFN3bcZf4Pe8yDrOAk1LnqPKh
JXl+1jwUfiRGM9Qb9Gq5yVhgMN1wIc+aHb6nPp5458IwTu4Lqno7De04j89rOfbJ
wncehApNrhDDToDufL6z9/f4F9wwgvaur7iNAgIAyZZexiW8+2PljUr6+jcKPRfT
BnxYnvo2MdqUr95eDxSmDSQw/oVrxa2qSBIAAy1oJSDm26c+p5K6W5PJJGe+zdH9
5MuopdVyMmed0jHwe4u4RXKBcqHIdLpzg8JdUSJgJG8bzf5ohHPGM6UHxRvgtGSI
TFnTSfB4NfyHbyDyA7Fd3ShUl4O5QAgevFBFFt8eoNyTLuxNYO+6IZV7f0mS58mx
8UdnmYq+WSWycc2MuiUAiXjtAprqtX0+Ij39pDpfjvFJLa3JlLHOS1V724oZ2cz2
Qv0rutOs92qmEi+kubnwiscFBot0n0msq/Td44AU3qV6fcVBqzyMyGpw4cJAMsIo
CfV/rrGGajdCnimQMwucb3fAQQsPK1ipHBqr4fWNN/50yv8BY7B8vfwVckYs6cQY
o/j3sjtB+0w5VnTf02MQG1h07kFK9zQK0HGNjGMAd395CgCPR3P97OqlT1fPcroF
xmfiFMC+hJFu4dduDBdiPbfijKgyNR6KwfPzJloYOco/6UV6WPUSncVNWXXCcJTj
0cLTgQSChwsrEmiqrYvGJZoQeDP+DVYy5dnxnJluG6RW7BPTnQZYyygl2rXUCLuk
5anbqVaxy2Rsje0XN+7FGAc+p8nFLn4asd6c06yldBc1QYwt9jF49VNO8p5Trzpl
JlTMrjYemqDohqyeVuZtbXGOpjnnCvgVHbv7jMOj06ON4oiK61pJO8odUwNgQWuS
vOuf3Tt+vxgfTfpEUPC8EOV9e6XBK3lF0oP1rKJnKIf/T1aQlPZ55UCXSAFMexVr
czbGKhsOwPT/dpcmsYAL75bt2guCjXkjPBjtcyTMp/GPIe86CGHSREbTrHjfemtW
15YK8hqmH/vgC3CVftY455MchqsTxJQ1ba8II7McH4PPVtxuNsaPJ7mCSSd27A7d
av59Qkk5cdhbO+B4aFlMexYT5H1NdSw8h8J7h2MMiGM+FvE2eseb4kE+njN0Jy8A
06EQdglKW+hypLn1sKnpMFYjebYMd67O6WwqNpDhylu5DmG2hqinASJQvE5g5Zb6
YB7f72MKWoZdkKJm8cZVqnynjBc3kcn07XzDrJIOH64w2NYsJ2fxzOVCsW4zsXH7
c6fye5xwe3iI50b+L2IJ+S+L2VepyrinUnN9gJfxqO9Czcp4uhzbd3AAJZI+shdL
ayE5kVIipxephuX7fyogw4Fi1m/hN+tESZZXtu41srfJZQbR91Xdp25lqCyqSchk
dYRwCMlWOuEUzaOmeweXgj4euagfdbxnVBWT+E/VHEYvp1ZflzOnWgbmVB5qSrNI
H9N4KVNBDyoQGN3SrREOr2nEJ4I02erFOGhIkUYO/+te36vlYeuq/GFbzwR78N6X
nUAwbdkmVz4tqi8yhCpFuvmOmicI7s2B2e5XyqeDXiCGizCKCLeShJQMin82zz0S
H5yKxDEk8gUfMfcXbm2h1loUbLqVJ0gP+9U2rEcbevHvX29cUFdUFHQbpFMKrgGL
0LotZdiYIwbS/TfDvbK1atjGEuoKsA/bOGbUovLEWqkdv4UjNnQcQDRGHj97MPzr
tRCHFvdMk+Rli/wwFYxePqZFvYQzw1Zw2Tz5KwlVt4QAqdWumUa/p4xkWUp3is3W
MnB7HJzjny7M2nrWaTkfAXIL3GZMZxq5ef4MGgMUOy9vhAL3KqNl71VlyMVDDvcG
bjrdEtoxqk00cOjLMPG5B4RzXnl8WWRXBbimfqlO0lDGy3QjDo1RU9N9FTwfyp7v
m12OvzCh+aYI1v6C/BU0mxWmiqZ4GY1Z/xJnkpNWU/4T9mmIst1YkdONA0kFxQ8U
3Bn4tnsib6HEnKOsg8/FK8PtMwkduLDmjhAmys+yKzEOeocf47kEi/2OOph6X+XA
nqiaJ6p1+HG9M6Szgvlyzd+StrwLacMvwxj/RNSL54p88FYIf1tb3LGnL2jKgaiM
u/hDcYW9ZGZLWpVS9bV2V8ectpbj0Kid8p19ziJ7Lyfs831RCHxZmFQK74UbnDCC
QACiHgT2G6lQzTqPb6Dzzm47s9K9qCL1bWF9xvlfIjZskiVNY5uj57zkSO/OuOdI
rStmj9R/2SnxpQksEp7/WlpCti86AC9t3ciF0mCi3DN/v0Ql71vtZ+LJx1+URen0
20feq19/z3gib1GF/oAFVSYPVRJgIIAYRpq1dqFRXQNGTqWUX5p/1jFHofItaByZ
MQ9sITLlFWJbBUP2VE39ejzZGk82N/B2zh9Ftsw9qUfCQnkcz2d8gJqZJpu+xWP8
pbyWrHBJs/nx3DuZUHUC7HWpawSd+tz6eCsOm9MEV7jFqjaPzyGOVmCvjI0jpTT0
lVtA0xTQAawqYP4nVQ4wKxUvhFmnieCMFx5lsQ3LsEkpkh8RCPLSUc6YUBce30dj
8+fdUprRIPLATOwtd6x6mX7xT5fcaLD+gDP7m7wDZWSWwVzzd2BzT8IFZ1e/2aKF
htyzc9Uw2whJO49B2S45UoAX31bYQvnaDzKIprQm9m8xRHgzWd0OzojlThUdA17h
e5v1i1WGu0IuFAVqCnz2I7pQ5zcaUthvPrMpLgYAbHro0D8biPMh1qfZUGiSL4g4
WOr09bJtRS8C9Sz9cf67ZKsCkcW6k9KNB96KJbnYiOwfU80olosRxEBng+SRyDFd
ou3hbOHWgzgrPAa+uJMIFO7YOE0ctquQQVHN3UxD48p0JM6dql1m0/uH4NjLWLQ0
cV9iF9ocbbWOWZK81U9DFemHta7HoDVOUqvy0eF0xH+RQwCaKmrza/TuzKvh4QdV
fcL0WHPRvpUHRaOZHliWEfAIZa/OkL1DFiPa4PjRMQUFvCOzYHJ44NrD1dfqHxM2
hE/4Rv2ySrDnTMJv2WQwFg6RQbo9R8mVbtL/UiP8l62RyzQ3brIv85Qs7B1pARXY
LDC2OrSSYPrE+gPh2MVAgq+UaqnKJ3S9n6sGVRag89b3t7ft7A8fpDN/bl+wK1zZ
Q0vex4HFCUrdht3WHTwuj7Ktadg5IR+RAdsyIahuhZqwV2BzFD7BFH0Px3Y75GMZ
yQklj5o/rsx/SkPTTSV6nIfVQqylzNj+nfzqf0Vx4lfxJ8kerb3aKU0fFtG+/T0K
FPWG8D4yqbuEIvAqB7kQpf41R2kEV1n8QWlywGPeBD5AdNoF1z99wCPU4kkcSHTq
W3joq+MMT7yKxDtMiES/MeB88WOvVCxcZK4q8xtgbJL9Q/rrL+P5xwgh/SBeK9kd
n3ZFuCHlvHvXeyB78YeCydOGcotAuSloP+NN6gKvCzDIqG2HjQ2zQF1F4ELcJtO4
ntp+G2fs0tcPUGQ8DAIhKLQ9nKh1WEAg2RoNyytKTOYgskIdBV2+1JC13IkMeABi
0df6ryvkOPp/DhA6U5znQhQRbIK3rzflBXV4aVc2XQYtEfmZCYczHhqp/uMymV4A
ta826gn/2QsQXcYB8WBpgeLnyeOHEoF4hIoLKmx3vK1pIH+oD9tANb1h0derc8GQ
RalEuoySc76hQO7RvBsCcTgl+nLkKGPyuea3Diu83cqtnDe1jN8yxN/1pgOuyMNt
paE03O6JDIn6NBLwnWPmx/vDc9qLp+wgYppYiRWMVOthw9PTSKUVDq/16/ANOhDC
ojwnJWEiErmFct8hq/+stxUCH9/W4mGoMZYNok/ie/6mWwOLCf/xwt/cVdfoXckn
sXjPWs/txX5IuOyFGBNUnxrLslfwrgwbxMw96z1M5UkhArrsjDSSL69r8r9ZYYUM
4uaLm57gCYi35HZhhei8Vgk42+xY0CRZjEG+BFv9YFMc80oUowFQpEX8HwNcU08u
j8zQ6RytLnQhBfeqBfo3yLDxuyI9g88Tdl3bjQRTcJRTxLqL01XvXX2THACTgXJP
hLzSFwvp1FetBXL+IU80QaLuUSiRIlkXkvIZ6NkxASXb5XgJ9I6V1392vfYDTGvN
yI8xnsGckG0sieUcJJmt//gcvKvv3UKwvMClSYrODx1Wps65CHvXUOQZKQ9GGeqw
3zOxdqUCoz+Y9zhMVvtiEFsafSLB+odLqoff0Qba3dnaqgsURTzbMoMXKpBTozkj
xmBLqIckfkoIDZfTr9tYQ5oA47M1T/1C+UwkK2eOJQ46mig9755y2dfEE3rIKdWr
Xtl4Z3WfHj/EC+oQTM+2AvOkD32tvIoLFdgthmSD1NJVsavNz74QG/P9hq9DGtHH
zOPqrlJN659t7xiogplMM7kkI3KP+E0CVEYpIZl9BMBLi3Ik+1EbKV1a9DJfxHpN
1ELwplwUQ2kMSu1Btcfnc83VwtnH+UmamxSnST10EQmJ4ea7yZwppDtivKDbjpUT
1IuAmXcI7xJWmc1bv1SAtle+FgAz5Id3JXQfrE1dgi2tq+O+QSgCtZ+UvebziBVE
eXtDPjakORbUWF/t65esXLKup4Qi0dQ1M4oXNqo9JqbpCpcnxoWP0RLolxw4go3p
3XWM8uPshChXh5gQwn7ae74vOKgbz/VrZ1gCNecrjv9M3FhFpHvWGJlGhWvzNds/
LOOaZT9XwZ2ffItMxCMIKOSXR7hAI/UXKvazzFlmaYSV5qPsgUaBU5sSJaqBeaOy
VRRCdiBCTXm+T7+NlPwPD0rIRH2BUdl/+i1V3wZaycbXea8zZHGtiFqtapX2XB5l
7+ytnui0MwKdoLK6bpN14LPTNDYRo6uzgu00lzBA272+oGNIbV7jGVXOGq/yNTvW
hJvvxHdov2v0DiZvqtJRKGsDKgcYmC6H+y+ziwksjlzX0aRVz4VVQoHrTUI/VIA+
8n2GOeRAqvvYxUc2kKmpGqNciAdbdTvTWBL5GyEyDLUTxQB7gSCg4AezzBRHru/J
kro8mNgSfpR6taO6j6u93afedk0/vGKcRESI4M2Enopwf0xTCOKrl9ThKowYdvRO
evX1hTT30B5gVZt77TaTZ6I2Ki+imnc9FvAsay9pWpw5P79mg/p8xXtxJ0QmogNI
koBgETF3Z8gIosX3bmCtUXnt1FfBM1J0hNu1hBwteP5tY/IlpO79k/u3rhzj/wMC
Luw3MjkOVPoTCWiPtDvVX6yv7lLrVihdU+hp5imtC5wkw8122yrV0RrlLBnQZJdb
TeF4F3F5MfVg4Hbj/QuO/flhdvYe+qXt5fsAE3g7X8aBSsAj0IbZrwTIaD6o0sZj
VU4YmXUkZ9sHEZ9SRSWpb0/woQq4vGPfLF0lw5bgX02CAaYDtA2iai9uL7AM6yLx
rCXVDZlkW/djU44sGOa3kU/Sdz2SLMFFL5DIxhJYuCCC9Lp/Q4JCcZZjmuUMf1u4
ceq45F3yVP5TGKzQ5PJ8LE6ETsnNHVndLaLHl6k9Dly6oDLbMtI6vBSe6E/rBaAJ
6AyeWh3Smz6TtQXUSY9Qc31iqYyRy0DwbA0q4sNmBs4OLOVmZUyeFb1V6YvVi2Eu
mLqfBht5OflkuE69sE/aB/bWgM1Q/Lzkb+B4YxtJseFfJWXkNv5G11giY5mI11Aa
63cYuxqHu/miO22j+/CVQr6zhQoUHrxFQm6FEg9zFYMjyHjzpDA0wwhGAj+hpsLG
SSmZ+I8BV8Hc9/ixJB6nMDskvKRSYjPFgmvSwbnfs6+HWWoD0K8Q2dmVpGfLb/I+
Rb9zKNpL8u7snnwYK2Xd795TBpGe7EsC+UPYwdfqpyJczdlSC4RvnSK4YXvqM8dr
PSQ00SpF5OooSnm4ylBx8ScI0mqH4UYr9RvQNh5J+D20bBOW4DZd9M4tY77B2uWL
EkXGlorymn1oZr75o2QmpWmS5BtKgl+R8f+hX2c6mgiURPBE6bKAM29Ldwzb/Wtr
3dHwdSvOUYsajbwfQ6A9ohPElnlpzORdjpsZgo1ZvonOecJAUUA5RFO2sXCtFULV
rrk7marhoHE6rZa649x/hD+Dny9WYJxq6l4neqhe7uhLwytPYdf0vqZLoIOndHG9
auU+V4EPEJsXDtXjzdo9gYoaqtK9xOWCNJRcqyGEFeuDSXqCScCJc+KcFu+0no/C
F/OFry6qw0lHqkXhrewnyk6PHC8iUQiVVtwLk+LypBupJYPMvvo+T7M7Uw1kjnAc
nVGHGsWXVAHcbuZVCkCD5jPas+BvZgzH4m+IWuFJKJWmyVpqtMIl3mKmTYxk+0oc
3aji3jm8bBTPGMxBdL88k+lZ9JIGg805L/pUHsZ94IQqndg6GWamQsFqi8yqrN75
X5rxs8iPWwOUZwyyudNnq/SZwXt20u3CXHPswlpZA1bCObW2xPGEiJL+G5D5WJEf
XPvQuBFf6cxoXR+d9kpkcdRawe/YEwkHT2dxm4OwFjaMnbjwwgyDt6/jX/S6bAYn
6HeEOe4L+dJPAaCJPOAe8ZHsVyn9CPljUDmboUpXp4hPg+6+OjX3o+qR9FoByGrE
g+iGvshFcG/Rv+mqUlot7cKxHOdkztiOR2pDG5zx7BcDLw7GRzBunqDOKK3HC6mu
5bQoIlAgBJitdSoteUOWF+sjQkxmiO6E70HjR6XcakE00De4O7XkEN/rpjxx0L/c
jKCxw7y4X/mvC4rkMqk2Ir5N3gfmZjtwzxBxu55/cGXjNScyUrr2EOrSjciNqT8e
Xtf+NKPyyfa4rP5JnqEVi0KG70CCBDHMRr5MBgl7VRt40ii8zNO6gw3IStHsjnzU
w/ab404MVYRGyl2i8rf4c6UmarVkkqusMj/mq6YwAplCug3whWw9ejNC+PTBlJNi
xif79/hNJ4YgCGEkvxYd5Zp77399bQdLiJbuc8hKN2A0iWHzfrBhaFe/f86MXzVA
Zo9OV0ZUdgCerM32X4YLm1spaOsOOBXlRwcmBy4LYhbklyzsrsj7yi5V4wT9gd7c
W/ycpy2G+qDhJu9QSTV9OcKbufMqiCOpFJ1dN0VWzfmHRhccqDK4eGkYf/ced8qW
qCw7/XnhKSq8XUfNNyGewXkx1svekjQxZ9Ch9sNGlQsH/IUrHlD96upu2VYffBPE
PnsC4Nou/SwZb/qzbEhU/9v0MyjsRd9RtrL2AsSC3yirhcvOGIbcAaF+o4MGCwe0
nDYs9mxGSDI+S1NT9XCsRwI50vmZAkiPfC0GZsfnbLBVrio2nVbeinDyEgihljJO
2OIKP6ZNRLcqkgGfjT3yKszY6YCEniAy8uD3xRsA/0mCoME1f0WulxDieu35M1s9
oqXK0Gb2MTYmFsCDgpd1RZ4uCp0gSwBd6Cur8jLNyPzOKusimHSAJu9wdBIMydpj
/BdMofFUisIzD3LZzIlZ9GLQd3yh2vNA1q7xdFBcfaN1X+JSUsosR60a4nIte0eR
WAjjOI6K7yAxKd8lVYmT1O76AgntiKl3VbIpwlRxYlUk+8OhbLU7V8sEXCcS1o36
fj8X33CNsQnt+3yADCbuKyzg6IxVPEO1ycQL7qBmLJ0Blm+SHatTQLPX4bv2mz18
MrlRu8OuG9CLqUIDciGZWmpHsZ5LGvFEZPOMJcJxwD6AvLTM6U3HuGUe62HRB6Qo
6iLjBuQIOReDdrKE2tOvSeKC7E936w+3yuQp8zR5n+vO6bd0DDafgUQEGFFvzAkt
LHB6ZIB5b41QPBTUOJn/eWVgjvx7Z409NEpntMbjK8FSqlYbKpxIvQqJLXJ6Kb1l
BOwIudiV9hB/XjgNQYZNLArbt7SW/kgXAgBFkgkSyaoDIKrZyyBqYPHgOEvXzb5/
yOJ/lLLUOWIUMDaYfWrJeNLl0gDBPO+skew7vqZzwA+x1UKhr+2DcdKT48LBV7BZ
cc3dQv/FVnIMtlm7AZ5ruP7+DrQvanGaqswQvDN+eBDE/+Gi61ShuoVxzMVTAa1e
ZzmmF3GcZIwH72xUO1plp0yMGhu9IiX+BNykUvqb/u8fT/XiMlQbsnya6TV6Dvbi
o5TR8ed7xnO15I73+6kcsjD8dl0qFDOsf/geGClkXAsjm/AQ9cML7MzDnNn0b2cv
LirLd98ucBWOtW0bQJF708fSAx3f38uz3ElUlku/PGjJEGkCOJEB5iYbqWL+ZqZk
2E8pPtVgw7RzPVvX1WUVYfYBmT9Y9X+s0vya/7jOR4YcBlNVY3/bFfdIssGXnhlR
5IR0XSQm7Ovw14PTNhu79oiXgnX0QcScLAviu889hTDOdm8qzrKQZo3eQBJXHGJJ
Y2BRXL0Z0DeqQPLUHXb/3q6wyivnKBBAx20G1LmnBL2/RJ9SRPAUMg1wJAfo3lNG
mThy0P8MP2aKO/2oHxVNGGJnS0o27LgiZi+Ln5+UKFu82bex1JR42ZLX3M32Bkrw
oL4bWU4Gga+jLle2wQDWmZ51HPN6iAq1yb3mm+n38b716Bbryr6ORRjE+KriEJP8
uSLF8Trc/AHAHh8Nd94jB9TZR5UFT3hVmuf2d0/BGg8hqxlZiOUyXki/v1LRd8FA
BszDjM9LQPgnpqflxJTUIrHtFR5x/lWaY2e5mrDN45mIJ4fx84OGra/Gos4NcMdL
HRbWcpM8nomA02DwC/m5qhTDuGroefqKBuCExTaZcX9EOPOEbxHNrWH04aRAZzR6
0g5a5mQlJXtK5HmCby9cL/gXR/qkjaxKyNA1GjWe5gs7JNURJQCJChQoXegXIs3G
xZ1ocORWNG0RX5qncQpsk0QSC27rOGNcQ9Wpxp1YVWfgyIG3Jtuxar4JSoTrm8ei
Lczl822Hv42PyW0A5bhUsqyyIxbb/QWT4fx/nf2+dTVwfWicb5EKXzGqnHaOqJPA
x9BJGy5Ehq/WKqlv0oCThEpCzBBy7uEv8pRNcjdTXYp/INeUV8MmSEjgKRC5n7lm
GzzS0JEAvMEiQpHyFevWGrYCto1ovld9xAEmAmIHDwNDTEc8TyjFXd3Pz5Ccnuap
1KFimdCSMapVIM4UCOA1yJN5TSKJTqAhdv2nhhAIt0//T6wBBVLacFcmxrT/3Er0
b4HMAK0EdCyHeQl2wTsFvk8NBrTROxec9jyvj+w3AHaoi+XeyR8gLPH3LCmXPr5I
ZsGKveWNUYFeTnWOdd5L7sGFAmCliBJZJmlMpzYteiY2IjDkgdmfIplht/uZU1O+
0frlx7oRoLvq8LxTEIzi9Fh3hE30dPqa7bfbgJ9bLw3Hv2a8a5bumZclVplDphuX
+leBOh9zipP3beub6rxUMd9c9+vVE49LMwC9lWVP023dOXqdV18tIyMcrzjIonV8
+IVCAdMMEZpqHWJ/pxiBc/i4porHIdr4otZhNgL0uMwl2qyEbUVpjxTv3JrKJAP5
4k9trgV4ENS0kFHZP0oVKNbaTcHLG3knOgW54UsGM3CyuHXKhCmz9CkHnaoEKjHi
lNlL+0zDRS9ZYRtqtxfdv2mZ1DsjDYh+tyMIubm/dfWJW/aN5+2+pls7e3ffm21u
4tZuSHiZdljFTien46dPOf7B/qQyg9uFE2yjzzNinzk6cVwJ+XteynMllI3TvBr4
TbO8QBtO5rT95exXAZaFTUo1cS2axGJkPbXNIK5q1Cjxdx123fPTZMXa/Jc0SzH5
FqOLBe1DWIm5FLwf9F7fcbR7G+NPj0vJZE3Zz+RwPpWu3jGnmP4yGhj212b8OAq7
xoshZQWhUALb1StDBaD0jbLiKs7u4L/RevujyY1dZ+vkqW9xpT9OKXe4zTP0zP26
2Y9gYw3PsMrF9oEjL//jPSeb1cRSNDTXIKskuedQFegIkV5jVQMSXpCXbFHIEgq8
eRZ3ZuNdg2opsAcRQvehqXYf8rCG6vVyBlw8JqvRaYRcV3yMDqUFagRstSR/RNEA
mXGtRt4UKAzBSJuicwjmaVq0lENQc6tYCdr4yd4ucHH5Lei9IY3f2NzCRWmVsKgI
E2WSxF/Fo7fWsaF3q2aip3bzZigG7gFi7WlD66OyxRopWPuAzeMle1CUipr3GTed
ey00VEbwrJi4kbWHsmgOvQeNQvmmmMevso/FDc+bcfFBS2bbNd5+FkwN4PwG+JBT
Rq74YEiO5c7iidiWocZdjwQU1jFrUdw/hTG3+ixSmEmcS9wVlmvkoyDtZ//HVfyp
w+43sT8HhBy2FasSw4sZureiuh/D/S20Hrgc07rBFpSkanibqAUJ6xWek+PTspF5
esknwA+Fhro5I9udE6oHUw5Da/EyDN3aiQ5WRZdME99zS3y+XGZVFD0kz7hIcRQi
QYhXTo9rUXuyWEaVW8VWLVZeVGtj+KlxfsQRE5JHCB/0xSZX2yHLETPCLqBJhtG/
bW+IooKDeCzhEI5rta27/dC4ZrJbr/yPJXv+qQNqdub1fX5Y4xeN14dy2dsAJelB
Rjnmnxo70mLT3jSkH3tkkIMkvxVhFGkrH325AxM4KMVi1ddqc33Gs+u+jPx99TTo
jXxk94uUNhPnFnWYY2Qt6Ls0H47BIZ/AnQWdXg1Hua3F5hu/M9J1QxmnI5+W3lac
Cjnm/LvIO1V+wMhUWv6faBOABTAr2kIT23AuwBGL8OxmDgT3kFgO/SrBr41OcHB/
G6V7aNMqjfLOPrSUzJiEYyNsRrDOh1+6fSnlbKzQRnt1i//9Hd6Pw8KywTFpGFtz
DjkuPfqUvIdr2zvbN3sEvL2oCuUHSLX4vFPfSLbpVWrkVHJt+R0I1veOSiU1XqkT
l7BhEkI9yS3cgA+WKnINtcbFR4u8Q1KCZ21+N9lHDD+cvM7qX0roTGzTpictY8SL
F5gzBT9qzTkHNW1leJ3r8MmGaaAh2xacgB2xGhnfxvaJrl+3b52M1QBi45hVYAF9
TNdEfJo580xq76wF+pVY4KJevtIsfFnLLRIfuI/nNISzKg7/7nFvAKpOY3Xja0co
N5rPdWs6ZfkBTZX+jWLxClTsT2gSKnUu5MIDIVQWTFJDSj07D8VNcZ3rUcD3a8jh
Vw7GqrpxP2jEat2fNRZ+SLFLTqQ6fcCqvtSMt4G0noK2GSGt+vpk31flgpb+FU+2
LoM8Xp//w1SSsI03xolILorudYx0DGBa71anvOXAWgv/BzClUGRXdUpxdc+frzBN
k88t2X+n2Wt9xa5Ol8g5bGEGxRo2a6KqeGFj+cI8L+KBtTWNv5CRr6YPjD2HVE1w
1BpHGlkyMZIBrRsEvfKW5DbO1JhL7DdYJxUq+oDD3PSZeBdlrdrMcHck0P9oF92f
LjkFkTWeSFvwbepYjEX72hNZ/c9jXGq52zvPKUBsqYcbvFvzcRm+q0XBOJ8IJbxG
/ffyKy4BJSuiQykBvQYjr/AW3/87CW0vzCD6ShzUIZlSf6BF3k7UhZxJEopHjchy
jkcXo0ifgMl7L7k4jZ5IcSngLj3L24kWq+Xt36tzNnIdNd37V1IiDPzZspcDADpQ
Q/gDIoRRl6KUN5fH+KGPIDkZWJCO8nG+snZ0bPcnaIApv+/potvvK1oz9AlDrIoe
Kt78T8yRLXqvn4MUU1NoATRb9xcNAS1O1oQUmeJBYXt8x1Knld6VvO55AmulXxGS
v+glgtF/IaXJRjJ39s4NvBC7iSV9Npght5qvl27kunh5SGlBfoEbxrOEZKdXQX6q
TEkFVGyQNn7oVWyCE9fpgzFWSyoVdCnU7tnp8XyGWi3a0JrV/DukrEGy5h1AU4EM
WyPU9Gu/yzzH9FoiDjcG9CxLio7mprzTskXR80QE8npi5Jql/RAeDo/yIgUIf5Zi
zFNJql24Q0IfrGUZ62Sn5rwbf3Ab2Th4t9If9Ex/DBBiyGlv8K+LAppQm12FWoMh
XYG2kCuGmjlTaaUc+XKQl69W6dRJ+QOhaxC1MJWSDCUBoablde3UGdCkD7azNCzO
xLgOTk6FM63mqbgRtDKLdXn6Zk57nwztHQvRCXLdWm9ruojN1Z9Ez8XHgqvCKCec
SghySF8ompm02Jk/y9GNGsE3Pvo/GdWF366jB/OLwuZG48J48RPQY/fEqeH1SQhv
L0EdqERK6iQoSLLY/6efE3oI5ZZppWjLuCZYoEYJfHvEXME1rYytJQmjobVPHZ1z
RhEDvKWtY1iOgviHGG9n+gSA5GeMqgUyasyxZW6Hkon/DYBZsBoF/lo7tCHOGikJ
9fj7ZXB7Sl6ik6+99El1tkELwFjC4dnMMCAaZen82mb+lTuWzwUfb2HOWj7ax9bm
kAMJ02qXNhSDcE0fKJybWg67hSrCLoSI8AMA6LPzGvvPHyXrCt2GoiTm8H0r0MSq
ozzU/H1mNgquC9Y155GOcMnpDIKPkugePNJhz25BnS/duqn7EF930sUoiWst+qfP
UyvQCuXVhtjSEftZfzKQLZ/LUZ3vE8aGOELEAL6Qw6oRjsF/71BamyxKdXByd/He
0Wc/EImhtoDOzpq/boi04gDODLuID5u25b8Xi4TpGUOqUEZs2MjOY6gSdKOlM8AH
2o7EVZ0fSqrreAqcism6vK1X8dL4NXFthy30M85apxityd+aARxEkY1r9et8NDSM
FpCAUL445nh1wAK1LynXWjxB4ibOF7G3XISr08vkWjGMgX3z1gEc/olrprz7pfYy
i3Ghjmc37udGhyfz+qbfq97b5ctdlJ3g0bIOH+8jYejn/qaKroiqqMWZM/9BgkE5
S2525G8gkTeNpwLuyQyhnq6AFiYp+6UILpTE+nTmBK+1HHiqKPpH5wLwYkrPJRWF
jUnBDooW0w2UX8IUiDVADYNyrfSnjaoCaLxUC0NOJPyYhoJv+BIl/MaNNajgc8fO
tJP7f15wBGS85AbCeMo9KEIDqLOfOuiSsUYh+VI7HZFX/pXTQZlNy4T6BXXT0p2+
AlyDCfasSDbDQyF/YDD4R9tiFLxqAlw23eVtBM9ZMn+n0FGpNs97LEchH95xNCZc
LX6Uh40O86X//eqpRSYYL4rX2FHJSBpu/JK3XXMAzZPJw2sljNXodL49ctBB+SzX
VVYr6LvdKZoM5Wm8HqZJ10quVsY8rVdU1BE1+dsJYGkHxbB+QJ5tHD21ylcDPSf9
SFXG94/WH3uKsEUvioULeejYMRwcNuVa0SSeafSgIrqkKLn/F4WO6tqBn29A2URM
yGCeTXx4ZcXfzY3vu/av7vdmB0SLBeoBrJrXYse57BCDGnJB46dByz5B9FcUSmfi
kivSX+HOnXc0PaQvR561M6ZGbMw4Q5Rgva6ld8NC9uhNpDfmr5DH/IIXxqCsoZ7K
P2zwcHViZV9Muq7wFjK2nafcN5Hbi+abGOrMVtsDKmnJCxsfU4t5wNeD5k/nfAvf
tCM1v2ZQo0Q3fStc0y+uD57ElCF4PQ9MBfbKL2ak8dzb+h6DEU14GMMH1QRy5LUT
e2QwF4ATasMGEEV8J+zKOGcbv9mF/DNDp0xbYe4PSN3jU5jTVtM2oFdqAKAqBnHT
RXwhdU8SyqxkpBaH3imVKjLWAcMDFwv2CsOmqqDlwtOubE+Kd+bAD9oNq9Ltsr2f
bGwPSz+dbX+WobPpdXmxt078dQgXDx63ZVrybAqr7oRiq+pm1lIqHIHtCBBoFm8o
YylHGPepENS+Pm11PEtx9JUPQfuvc6gybed0PX+h1WT20U+2bEriBlFUeGARqcuj
3eJk7yOZ71TDrd2YCj5Vvj+AgkaHUmIeuHlOFuwN8d7xtItY0DG5PEa0egd5oUf7
tZHfsBHJmjLGlLzSlAqNeqXYQX6ZAVs15feEWdTLT9TsnEcSHOcg7f4ivMAkYGA3
YZhmnAHnl/+tAoVtQu6WDfQGw6W7PBqV/2vQ7YOAZB4E1WbsDx10xTgriJJPcjcJ
rx2P36ju/FjU3AnreVeEW48KlDfPyD6Qtco8cKZRukYBvB8laSksSIa/X7Un4ti+
Mxv6p1fgo9EP6hNkJU0c2e5RZPqCLcttp2ppXLmXfk1mMkkw162bNfWFhwYtiqsP
VwzfXDyVi64h7abtc9mgmXDFPPgKg0x0h8nnvjNri+Qmt8taG77D/G8sDAYEQaK7
KZoM0HHmt5oWwFeM94JJDJmTLiWSZ1rDbomjmliujPZVVTC3YQAabfwQoMOg10PE
7GBSeMl9Zt6fRaDzL0bQDxz65JQjL2UMGV5Vdk16Qm9MEvt/lpnDHr9mefUwMoJh
177E2M9RQRGmD+xigpwMCYUDMDcXfpsoOIfDBxe9I1Pjj8KLa95hf3WtIR+B0Dif
na0l8lfB4mVy3fK1WqTbVY+Ih1GoGC3RgD0Uq0eSMHBGt2FC4pCia6J6ZOGnwnJF
vUvxxnIxCUtYUIV8T2roaPt7aNL5crVEU7BUgAdk2G3idpTp5JTjbi9mgd3DWl8+
nID1x4TZ/nGIfTVoqVqUx4rcAUXB5lSdlmQmpD7/53LT82Z2ESu+oRCNJoKxHDkz
1GggONo2vrtjNmlgcd2IvKlDGmpopVMn9jYuRO1qZp3HQ3nvTLCpp/m1O82YwFhG
SORLFj5ZZSXAZ0qWMc/hTnCl1cxR9u+VmdJLJ+A0uAcsph2Sltd1dPGlm+J4Vqna
zNU8ryMRJ2xiH0mH5BXRhhLVYDVSYQQuDehr4Q72t4/xBIEDPkp2dUkycLzj5Gek
5B4tDAgrwcggvSzD0F+fg02VduIPN8+2frOgq9iJPA+URypygy2xojzb4yuj12ni
4MCgI33l89+4RCGhNPWoQv51yTJooAyKYxHyZ19hCw46QfBO2FaAlTynfsAwBfvn
R2qjyIuJKFKmCGx6hbX88EFIVPPwM7XIqcP7OC3xPujcd+bVrk5PviEBt1KpILMN
AlCHqZi2gXQmVxjiZDk5Mjk1P4At3etzhYGNFT86v1YLH5HCZgNCr//2zU9ylIIs
Jwql6lNcNgwC6aQGcF/Gw858bSHJCn88NT2CDTk7qvpBr00gqOZ+vN8iOmE6uuhc
cMRKknAMZizPqoU9Zz3hW1bGiuhkeRZyHQOZ8Zd9LWRXTtBpgQ9Hj+6MUaTamsS5
EzymskbqDudGwfdrU2iiProrUMfnrtJWwiEcNzoSyqBD/9syQ/OWwXgC56kDuQsX
E1gmvWKkO+YNigGBwT33dOEEkEzFJJmID/XxyoY4tcMY5ejFNioeCwC1gU8pT4kS
dfaiX0/Bx+EYAVl7EsFJjDCWhuSpuEFiHU/9fgM/ZME3u2EbabPSR9/l8up2SJqz
luXZuKFkfqqq95ruL9G37ZL1OriGk0u8Yzf7XWC5+ndtWkFISyEva7z66ZCH0pMC
DdzlG51nfVFrR0xYc7sr4Yfrtakh3m4W+raKml8mRrd/oRpaZhwzCnjTq2HEYKil
1aYMzvvgUgU7xD2kLNtwoiDq50IlRYPjFnk5uX3xalYpWQlID1Yy6KE/RO8uSY7n
euScKtVSQriAxej2s1/WF1QubWafIYP+rwWBqi73MvrJpaFr81mXT24zg+YYZTeN
QkgGP8gUncp34rCL1rrQhrSj5MKvbJ173wXk8IoRlMwyxRi97ut/PnoHJyrI6/FD
WxGBHvnQcm3yEG7b2UT/a/pDvceW49uKiDEOPlgPcROzxf/xSRpCMW+aTwxGpqRw
6YbvzdbH9wP2gnJjS8OVR2TM3tET19qjoNaqF0uyyfohdPcc3Ggqod6Vgi1KwI/Y
1Z/C9Z6k5lVvbfJopaoqBNwnKFL6Ri+UUF9bfWKYmAl0+XtF5M2w9Unu0iRxFqfR
5DpmjG8026m1nRq6O2PXINZ1OicO+AALtQAyh63Axb/6ipUou+cUk4pQH6l9a8GD
MImYk68ahKwfV3xzEuaPImEl5b3E5aJkHxL8qevCXko3CXa/T5h+L4KjmLw4EMSk
hiZ/gciPnYc4TxxfKJG206i05tAUz7M6thvW4SehN5bIL5Cdq5QaIYzOvEJtnDse
dbB6gS6Z9tKqnBKLPGKXeSQz5EJb9zngkvqHbCNpbwPd0Zcj30UrUhr9qtXOE5An
yel3qgGVeknOBEX4NP51pzGuwe92qq+UJ/6+3TeGnifbElFkEGuKJsCWbqqa+YJ6
lDSPgpUofMQPqz/I5PLBf08uG+Y26BbYVqXWthSQx/em+PuRP46igF0oWjVru2EI
v7MkJLvDKzF3q51Q0yKYWquaKYK2vRgYdh+OArsFS2LUXJ8TrXU+yMwjdwUdbtqy
1zDU4RG/kmC673+YZAWt1ELgUEyUuWbKmPej1nMKZuG7NazP9FTGTj1/NoG1rBpN
S1FtebCq7DlJgy1EiYwI5npOePAmwVdW1TghvUokP9MAjqNA8VFakii6sF5fl8mR
tKkAR5PecwYjXKtxFvt6a+s+xGxbWZf9NGG/V1TmzdMTLJrEiPjg6PfIEC76yyWc
1UjrDNsBriY9TBoOXwCd+2Plol59NE7NmK7X8crwX6cXurouUN3RrGmqLyBFDNhl
rDZRvRHhUXnFSY5GTKKrRFHxC3WPY74MmE4KzhalfWNNAqjBewV+iyEsVVhwZ5/i
Rxi98iQoK6zNoO8rzvdMG5yMTR6Wm+14jTnVKeNuFvqT4IjhHhfOCGdXAmakxKsi
3Mhk8JhZyT5po+Eet32v+sebm+tNnrkvoOZ7jfXN5LeSwq2wnFmyR9NMCwSYtB0v
2qtdT1d23EIaYPe/bKQMvK5dPW95wTT9m3f7MmVGTvOWCO/Z5t7zRZNkz10thQZa
O+gWv6nTyS69IxQ0FO9LZXksYAW69bWdiuvi+HG9+Y8h4zQOgY6O4JgA1U69Zs8s
a1abr7oYsyRrJo9koMWu+lY0Wr8gGXxcMnZVpxiApLLuNgYmV9IGwR1tl9lfQUY7
Y0uEsS8qbxGKQtykVzs+NxJb2RJWtVvGUn/HTBnY40lOT+AltoQ/0NFHYmFWkPO3
ZplT+jtcU5qAGCgjZeVN2IKpcYiMVFfznsGi/85kkF/N+lBAbwP6WNLRYOGnsZsY
vbfDAWWfn1AzydHnZrMMKsPmIKk0gblDY+158vSnVq5hpugJHfJOE70OKou9c+BD
Ezr8cd9MfdMo5BcAzR63/+gd8zXr8gBbKXpaaTIEHrCU5EO/vzpfakFYkmaqx7+M
00w5hl9Z+l+obUp6YMzDj/dytljY+HtB/bMFTEyZKwxMRccz0aDj6HLJRNMyDT/U
3nKOPWRpLdxL85bKfL1YqBdmf1lfEFvTkRCpA5gagg9etAYpRjkUtDr9g0bB3h4/
ZjF+dt61hzcBe6TWlXEx5zrVgR86tdTUmfAtNuJebtc7N4GSg1vWPbaukb2nvQtw
zytuqTYRpbINM7YmyBzFNyC9hzEStiTa6Zts2zoUAj8Jsw5bC15467IcOGRoDSej
hub9wcp80/3vTYgst7Nz5GLj08x07x1vTYyKw5VSVksqdaWHUEcayjZJ5U58jYSo
ZfQITuZmCNQlI+8pkbaZGhgzcQUnZyEbIH3LaOLtneFNzR4GdfmUocYnvD3CgGWF
0Go5m0Nu+iKY5CcB/mA/iNo9Q2CSv2vRmwSSzBFYiWVzHCmCHlW5UPIq4I13J/E0
qyo+DOLT4QW7haG5jLaR2eBouuZCEOQLesT3JElCFWq8zNSWRdi/fE+pZavfsbII
KpwLETdxbwV2pQDIFbTDyDUsqqUMk5WdaSpMp4WtLYeNTEQ7+2WnYJbOmltUnobq
5V7ad3LFoc4JL9P5KVKhUIzUOkFE/wTjgtB8+4oh19QrZKIuL5mkMsF8NO58+bzb
864eEGLqFrqyqvuSf+RliIZ9jn3XRyikM2OogCREUwGjyekPS3sYJqbYWm359EiH
MznwhXCU8KDbnHes82m9x1zzFSjbMkK1cDopxWbRoiqZqi/vjLjpvStS8umjC+EF
3yYRy7NYuxfpgj5e526eqehMQmiXoqgjyIRaZSowisa5mRQp0s3rTfhFw++Ul+1E
yyhJwij/eljUj6xbjiS8IAK7wNF3/lR2vlC8huUKq3ky6lGWPbQbOxiUf0oWokUJ
2m0vacmm7Kayb9WyxZiMeWWqKx3ZJeRRRdV0Ubjailf9A1ZKt+eat6En7txLYxVN
DlwsINd5TqeofxtFMWfpMr30B4oWGoR3YPb2g9qspnwA/AFR4QZ2jjGLyoM3nW+s
uIVkgpu1RifJtHfGw9rhlvd2CRxu6ySUvSG8rjYE8A7s5vdlwxPhsXIDW3a3R+K5
AFXoMCCrj7w5w343L09z3TMps95shYHhmebi8ZT9CUA5uIlVffN7ZOn4dx5/HoDe
rpqMEtw3tVHl+glNsJ6QJPDTAf32cnEcc1PugKpQw5BcwFUWVluceVyD5UzS0t0k
pb/JKFOmhs14B8gguQUN7xPa1BHWLFhFGNExZ11jVafzKHwmDgny6i9Ddp29fRuF
6kkXODh45AbpxdZyxtct7fOb0IvVPvZ5OJXU1HE5aa7dk0iXvdEqseLfPRD0QwyY
yV/EoqppspZpWG9d7bzI1zfPL1ewQnHRSwMl3s9DiFzp5uqrQ4lbEpYslyBbSldV
j8ZK4/rXhW5QBDnBxyU03Ara402z92jvvWyCgnVMtxEq3Q33Yt5hHPHKHmQEG9Zj
KtsQmgJtSn9KwgPhXKCLprx7KSide7+xZlw/W3fsb5zVeo484RmeLATj0yb9+F77
3krT27dyysSQ/S/jdZAft+gTwOBAtYhg1VKemu/CqpJhW8gmOwr3lhD1rdpBchBi
PQZ9aSg7hrLlsic1RS3mjtkKAXsdfhprz9uIFB//8WXgroXffro/rQjF9qCT2OiU
YTbi5qt8gZEZVtOK0+XzJ6rzdunPgPcCZobVMlOMBKq/evQZi7zoP1IeQgUQifLr
5pkIE/ojnXKlgqFa2gxj1MogLPnKg8KnHT4tqI+sVAiezRUCFxS5fJ71V4SAJsU8
PRrx02vfqxmGRvMkCiwBoKTPBZKvPoZEte+53yByee7aTdKLCBPdFuOP2k1d36h4
RaKd0CMX5/0YOVCsEInCm+SWs410IikWqnGRwTkTbvQxA8kVCeE8lPNwhROAXlEG
Vb2gN+tHMN61R9SHIMMcN9SmFl2Wr2KwJnHMJvEpg79wUkptgmkSClsvrs0lezDN
MIM8+d00LKZHXggUhR5ZRqOxdpmrjhUB+Q8Gep34ztBq1UxZ4toWuB17Pgq8KqEc
IBckdS5nMrmCCHbnYRo6oTg6dP14zo+xFQ1PwA8hEouJXvltGX1DszQv40eycvfv
nUDfW5uA4s+5NRORqUx6UEXpW9ze9yNutmJ6a1C0JU4+AQmrmwJVm+Lg2Z2eWVcM
BjtPcugDfw2vN0f2Q9DW+TCaVLYjOXaeFvUDuDSsSAUdeY7/ezkZzl+dYAT/6vWW
nxKbUH+V/JPtoeRWIW9/obd8GEbET48kZLNnc3ro6j0vExntUuPBsHY/EQ8rt478
+sfKi+Hmg2hlqvY61drojrxLGejDi8XYGG0wo3JZl+blEUYTME2FmMJ1X47t1fFl
G9S5wvb8Z8MhBa3q9ZyzpkPrOh6FZl4+iauCAdAObkVfSrsQqcP6JCRenQbAKbdq
yr+ILlwVoglmsRKIWNX8biNxkpAboWRvik+f3n/uMMrbJfJcwCCOU+275TOFGu14
MZdamIRZVrTX0chSfuFWQbAiodlMDVE9ZdAZsYvGzveKIF+mjmTxrm3lGX6du244
WcLbIsrLqi9EqFS3/yyHiYklJBixiiLMH58dC9riHsa7zLnCBG7phfZxiuorf3jl
O4cqvuhGsq34LuBrPm0JMRNCY0P1w+oQlDXOJt8Cvfd39DOawp9z+hMTNCgKpJ08
5EMoYLf5/SUkUSrOLVJOejrQICmyX7fYHlMkZwycKh/bgQitmRVcrgtB48t+mC3+
jZ205bUq7HwDcMQUgv6IjmDg5ydapuqKoPi/fuFRJMST1sn9cDMcdjQsrzWeu5dc
BPm3dq24DFsHbztw/jQjZmFbPdZf7NilQDu3Mliuon/4tDzRczFiBWvfddMdkRxB
EWOk6sbO6VYPe/Jj31+CsSsW5vJNQLIJT6B4Sbz50MTWHAmMRt+HMTjr8XiBGBFU
xYptuid7y9i+D46fQq7ArdsJaCHjN/GT2mxl4MbjKY4hExNiztWXclVFBriyFOg7
WCe4VEdxSQ1eZHwIB8cG4WCXGG5lgwFhonvTZpCRSQX4ieQ05nig8WthEfjJzh6h
Ct76T3IpiOamFmGgBzpzB8Hd5nHaCz7I0TAXZrDb0rPQWeU7+cePiJG7e2pKkSX0
G4EyuiGVpvj4VCwasWQLuUxhW552apSaZjDB0KdV+sY1ZGKO1BgUcaLAKPCfbhuu
oI9eC4GzHIaYjjdZ1HU+R7zqQsyiiCjm2YLPbRBgi8JOUJ3MsJXSWAJz7fCMfoYt
htrpVc7Hfzfe2HsL7hbnH6x/MJjvi1oi7wsaL1KxH0/iM1ejMJT/5NtQhnt6Zxp4
JdSDnme+P1x9se3lyul8BcUfZ1vngrdQPJzxisjRClp0qiXbQiZnHCPD985X/rJ9
kpWIW5iF2riUTMnI/w86I+EPEe8gFIwG8kp/ctKQIujmOJZMUKwF4eGonQEZgo+Z
HCGOTjtMVWcVFUiLAlDXSobkiXSUhxSxdiNmXPrPe9bpKDR3QuA+Ep4amId7HPjF
sUjS1vhpnNVAwHyPZ82ZQKfHjmo4WC5iKL5n7kpfuT4P3pRSFfZtYTiY9wP6++K/
yHWOFBuoj89fwKHY/0OOTBykjdGzZH6+E+/42GSxZVEMtMXOYaiWLERbrlA8T1LV
5lsfO4TG0lnaIjSZB54ssPNOEYCli+wwRPK8OU3yvv9xxk3VaeqkxzqIPSrqD1j1
4tGsO/Om7iLw7NtU3DqRCaDSGJDHa1jRg94ryBNe4WdffL67W96w188IQjBnJhyK
fTNRIAAcjSdqHlOobHqK59vIziVMaIaQ8BDftL/Ql3gKGq+tJQaNGi0yHaOAce2z
YN0/1AjO/Wo+DRSRLxplk2m7YJ/oMC+Y/dRQvE+6KWzoXs95ffiUcS70N4ecvhP5
Zp5Ze8CBOPh2ObYCKOShikkBbCNmwMGRGWZKlsmjOxBPRh9sdkKDPYnu3qHLPuqu
nOiHYQ99qHak8q5pIw3ZRJv+Bn5XMHy0Q4/yDPkQyYj24ajib7mbUl397gYeJUaw
+kZG6yGeTOyVeCfYKn28ut5bmXJTsmyhCSyXo1a5SsUUIeyjah+F2q3oQGcpbQ7q
Q02too19x9gscsIfSu/0pjTrzx0SYGD/UCmYh9SOQLhIlJ7MmYgbZbErgekBp1xM
99z0WhYtNYBoiGNcMruRsiqd0vSU6G52/aAdEtUrTHSOqT8JmO3qkTtldx4jCyzf
FxOdsVAQv25VpyZHGhF7vSAbw5YgtEBHgf8Eo71f4OI5Uhl72gg6yQwZpXsiQq8H
UN60l5N1miWTK/CVj1N2VP5hKnNsoOmnnexbWyXSlNoFtusahPTWDbeksgF041cg
OtHyytcYA4P6ko1M0zLMi/SUoOUvYgA2zo+/wV+LMAxJl8OuHETL+LceEVS1jJKP
+HluzDeXRnyya612Ox2P6uashGb5AVpE/ETwN588nQztiyhMhHmvi5YT3I9ET40/
d+KWVX4X7CdxYFlAs4+7x5HkMzYpLTkc2e1wMCAxB+Yrd6NBYlghV+cxURKWGZzQ
Wem20zLnFYHlzbY6C16RmUE5GCmM2BOI2r9qLmyRCwHFna16QnfxiYyhSQV9QT0M
m4aul/LqIKU7g63TI73V03yyqXPK8PpC39GW1t51bCWXCSf/vwjOgecOhPacTcNf
9CVxKpKwhXy0lbQjfHvmpHlelYFHT61e6IM2+cfBC56NmDKe39R5wYl9mDEIgr2y
tipvzRCI2rQ/q7R2mqid0A11rvX3fQXgdek4521iJZqTUWFlT1pfuz4wTY/ql0Ha
tdCfx5JfOTU6fhcDZ29ggI1J9z8zh3OJW0kivXDVoQk2jajMIcCXsiQPdzmZq/V/
W7P2IDz6uRv+CvQ6DpJ96QuZ2sTw79SoRSFSznYhq7Nmiu/xmde3nUg1qTtRfcLU
iPR4djMRjwp7EjZPM5VdNgCRLA6ZUdS2qc2evupO6RmoXAFXtKHVj2VPnEp24GEl
c74jwMFfEZyPDSO6kboMj975uG5gjjYU6n+Z+XaXgBb5BKLFAMzCp9dS4ZbBZ6XW
RXhyU6xY3BhAmMWpa6T5MB7Riz/v5539H5TUg4D/dOdDdMy6o1IajRLIu2jUDZT3
VA2szsgxsm5IxT4z78RHG/TyXj5GqJ9HZtBKamhn3faG5Aay5Cwd8uR707cJdJ6F
lR4sTXL+MYoMvBUFNA4539BFyCb/m8XDfouncmClzs1oyNdhry9yYwUrTR/ErRFf
zhlUb7UUPejTOfCeRXcArzPswFIM3DgEKfZLYqmmKnV9CVsgqrjn+cGp88rSftuK
3r+7VoRYp2VwHo3JFFUyYrQfpEkyhclBce9pVDKeVYsZkzupq1XZPeVNgY8uIlmZ
t5sBRS8O4jzpwh1pGuMSJwqX3U5pzRFhT/3/CsXn4TbXui57qipP/DpMBY2zw7v3
OC3Su4pd7xXhSnck1Xaorqv2qltyyvFQxSdzJDvQSmxU3PO2/DU1GV0bChVRxBAc
JP2MOW9Wr1xQjr01BJwp0MuzPlek4HM53te407rW4XvaMAI//OKF0HjX4gBuSS9E
VVzQIMF4a9t3xttF5pT8NJyZ9MvMwaXiDM90TFMDmvp/QcYgqsszq/H7gQS0Qj+R
4AGTEKGIf+RI2wtUFicbFFGmEvGkgN3XSOA154eomLUsPbKPOekxlFu9l9eTE6yF
W+uWPhqQa3rjO8kdF+cBj81tAFabguDWNZQb5+/8/yBIsearO3Xil3Q50+72j3qZ
Gwi01/sbPfIW4Mcbbjk9hDeIWQ0q3dwerT2HONfK3ZVnMjHb0ACmd76VENYGQPzM
7Nqczt0VAq61cfz4AcELlY5my031cmMqAoXk0R7qvflOUpDvhqhudNRi2V81aVNB
wvciiHlK1OI9bZwqQFQC45DsEpNaH6T/gpEdrKDbkzeqwFcNB9dS1MPbs3jOPA63
qHIg+hgf9MVPu2TWKSolgWUFmqZ0Jku7gnNrqwO+GRfEEmiWsOPSggxXWct1rDI7
GPE1n2TzJR3sJuqcLVuDnWGF7SlgP8c76/dFyugJ0Yzrh81GLamJkcwug93ILemN
gLpgIwM7dk/AY34ceL6bmkllcyLaLwqjDokiY+CsShExN3a9j/PMWMwFLbr6dqy0
PuIci+Q8VRfBE+vFyndoOrISDkKcTS3LLEYMi4bEV7l6guG1H6fXtgCSeydH7r1M
ceJLBhij9flbWeknOSOlcsYy/z6lEwYWVAClEEx2akMy9iqaNRg+a0Je9HjX0tvp
rFc0YSjW0EuTv+UbSNW5b27zKUaPztufpx/wDX9suCHm6X7TnSbpcEOYB/z4jxYA
5VvwWJiBWz1jNFcaWyKSsSCwV4v5/tSDyFUpUre3RJNXlA8Ksj1XZj58YmzEV80P
8I0aJu95U7+HQbI+81yZG+j4g8CUnrwnjGMPBZ1jp8hZQGKOUgfIyD08ko4BNu21
IIF9qpj+HWay7COVKnDnPysgc9hnKtXlEFNFuD6my+8GVwgcoMo+7A1Fo8ZTFdKj
Q48f/q5TxG18i4vTFixSp286T8aS+cxN+oz+OXGncqQTGUmJynUMweOPbFohmzVP
rt1wVhj/5wHbZ6OG618WKBVHVR0XpRTuPdmgG0QVHNYSIJb9I+yHBkmAKKebBnj/
nh388v8PI1YIHeTFjqb/59ayBPaO6Lf+0F8i+cImSnOpOTyoNTAvF7wColY94f1Y
m+LqkS0OfeXPjljnc2VM+CQudml2ca2nIJZ3tU5VxhQ4p6+ub13Iz75LnGePkDXp
fBrJttZC34rjx1GZ5uJEHueS2nrdbeshBXngc3sh/vHTsagG3p6j1nlXWTfLW2lk
59b/FpqkOq+g0iRMGa2ey2WE8fnmeesbI1GIDcQmF2k6R739FNLeWndk0oLsqoDi
0rk9/ytCTvKZZiXSVBshtZiq4ZX7PlbFxmaWHYnT/ChaISb3h+jPQMbSiH0ZQFN+
W4tPjQxgiodFLoGRWopqspNOymEIcvRrA61aSiQIkSOZcVDdnr98FxA3d1+miF9o
Fgi7YvCUANz0Q3pT+9Cya80yd2OnhKeR5H2MiEiyJgJs14bLKcBNSXDe31Y5QNXP
s13rhJ1omFy40jk0vnWjRIxl9QYmOT+5bcYSKYQdJsuuP2mbG97j1ZphvrSboBK0
Uird8+GELfrmsRhioz2htaCPhBB3BmOZFGISFo+akvFFBs0OnUOnZymMa73ECsLm
8ppi0SBQAw/Hgfat4QyIVOkIyFsVJPAiOWkpZRhQwA3uM9LdoMUcp2aukIWALyyR
lPSok8RBBsWDvp1I6ZXT2fS/LprRpWPXfcf3ahKp12+zBKKwgEgNi7UMLX/k0TAY
q7pLxxNKmx4GtCbMIzgjZ4MFZboHHKID4lNV3sR9uhTizuUAyhE1FG3EvDW3HgVi
rHMjuUxSqx8UUMnKCvh5OUhDVwNTGLAPuJm4vDCwGbb7XHe7EKJdVtEdy8WMOHfH
9dTth7cPTHutVXENAlD0BmEQOsteRi7BY1U5OMYCy9e1svKwBwFl3il671X/Qv7k
eQubd8f2MHi+RRtUU6mslSU/fOp6FAmXO2hDXdM+kpw5BiQdaJQvQhEkol2Kyc9f
A9Dt2HY6MK38MMDFnp0rfcZAY11r4dJcoN2ZCbRFkcSdO1CAE01rpUawFOnx2VO9
LenDrspcrGJ7NHCmuNjW+d2t7dMeGZdRAp9SmWU9rec3YFpDk8yCi9GCtPKMxQym
Mjp7FOXxXvNP6Am7Q4wIBs7div81GOqlF6c4ZNWOewA6sf6PgcT+7UJblgaGLZE9
zxEcPxBkFpMDHluog8UyooMWpVVGYNathA38FucfQF61BP9dEuymNoAebtFTkIUL
zzFst+NVzltchcg78W9MLFgchvtUwQOf69S6wH6iCMcz1EZw51LlYCcrQ7VLIGF2
KkCD+/zD/pqBRDNZ8/RZ0hnrl7smB88O3GXJWBc7DzFv8zAc2NzlBEAKuX2HtZs9
5VsctH+swq/FMUMZ5bR2F6cav4dzFAgGfNeAI/vbvmgOMnDzi0jGyhhlciVaDHpu
ZQu+TTOYHa6mqE4oGn1Fdqp3GC3HCoGrjkeBAJwj1Pp8aYyRUlMnv396XkJvrAeo
BuXM8pobZjjc9zlBgdULCFwFgm2pi57fVWN6Pbt2OUtYBWXFGmd/LWuJfAPVp/gT
TzH7FX2YAXbs4yNvoVDx2AH+SNdiIcIdEaCy08/Y9PMHQtzSfGYTixgAzGoxc5/t
DOZRITLd1Pdg/aMjCnb8Ouwzyed8tTe0zJRikbngZXHsUGa2jtK5vuvkb/A/TirY
Q5MUrXmtx8fjRXgKT9s1kHKe4KFVr0aL9XvMT34hYiT7H2urwLAq9ZGAiYXUTYgS
KU0nvR+mJZApyQOaUq6jwT1VvCZf3kXANJcgPGUqtR9L0HOTuj9OaGGL2cK4oM3h
UST8AAjRGjVDglM2pIOAhPlFAjxLIaXtQcDjhd69GjI4+vrqcmQImUFB4WcIUm/s
mX8svrqz+yKEB5molDE/SCE8VqkEfqOwhlvMpixr8aU2ExlEzPdty8esNpFwitKi
IkYkoF68ysm9XJ1632UijuWv+/3aa7mvMVuGFm41xLCKo9YH7Sr+GP/a+m2j4zej
BcQG00R5nNmaOrgtJ01vOGzTCE0bgdQ+JOje5FdTvqy7IBHka8CfMzLFYzbH3s29
bOemVC8Iog9QfxR9Tfex2uT/OPv2AN81GfnjGzH8gEA9eS+CiMrp647FosJSm5x8
cM/YK2cNI7meJwabA81fVrfR1gnQaEXdRr2WwLaJEBlHK1mBye87g8+bEzN+LCWD
CfcomU8fNYiBb1VsBb+8hDR+jqBnlGC513Ojr5PpOoysDpmMBgQpaZfd3kyS2rhI
DnRwfYByiQg6urDYiCgDZVX9Z8rdmHHnCIxEHvVym8JgP2X64t6ASEgd2CH+1sUx
bh5YNOI5ZqEYNDcQa7U1mWp7gDijdpwADm9JZWfoioR/jllIezKKGsIQsMWXrQGx
e61WoP6QfSrzOTIIq3pcFKTS+Ys25QhoeNPuhkaX3E7Is2vQsii3N47+cMpKw/X1
U3QweWTwfb6lIbyPBliIp7kjae37lLlMSqcha7xRWBb1CGEva1/tcMsQrF1QNdQ+
psZ/J35AK2omsHtwYH5kU+7bhAVB/MCy9JTlQoXI+Ape5nYd1PupQIWSQq0zQw6p
9iPmHc2DyjAX1ZIERBM7EcOEgCUZUJF20hWBmqX/xr3+cR03QtzPy/oKfsmXUKXk
gisZ62Mt/zgMahfgJS1ldQ6nx772t0dSGpDi/i7MdDpzcZ7Dd6cWaURfRQola5+U
fJjhJwhb/DCpt6gIeIC/c3+eMERPtoMNEGZl3M0M0KketUcuiVzRa/hGAjtupdSn
0b9atnoJiK/qTozSYU4EyA9mPd1/xwToeNjeCMctZdLjT0wqxzqyWpDrbAS5HYlc
9QzIDldj5wiOIr9dMDKZNvRH4ehcJT7R0RUVnTZ8lvy5M/H06DmI4ek/FU+RejqQ
+UdZVPRULEqTvOAxrfWRE60JSvGsPY+JHIISoafI3qwK4AUAe6m++hI2ZRzGflzW
4ZJedB7V9FjAozU7pqvq0VCrXbKUENeSF0XlF7d1RURJtim1seGDSZ5WY2I0se0p
luboopqIcDmXvp/OtwahRg8DogzQ3wVBNT/lNOI+G2dcm1OveD45Ur3ddIy8vVOm
9fL83JF8OoClNWh8PUdMdgojQOcVC6b5Xo7HKl0vNVnJZdltrhr/RZMhEXfuQZtC
8QzOZ0rvaMSSNLYHW+8DfBeBtW7PXGGvCAnAtVjKlDLJvuZCEQUYkdPRkpoVOO5f
aYuW1/xhl5UVTugt+THs/+lTwk5AG9l0iCND+0oa5rR/al5URAOsZM04+y2VYGAr
NsQNyT7V9USB5lyK6YxIREgT/YyxHx2D3hcNIxgiK1HzLf3a3Ke/j3smo+Ru7cCv
3W51Pz0HbTZmGzGb30QIbKSqtWGa4R+0vR+dmu62Iyw4Mz5h6wzSOqgN7VDzick0
Qdy2DLlRjUjafdQJG++PmKk3Z1avsYK3aapWoEqs/tXB8K9G2NVc8aFAipguC4mJ
xs0b3KreVgpzBKFf7kZVGrxiJhUwfHshwf4BtyiPe6JKz9QOwbqsX+XwzC/q49O1
prcDoZl+H+DUpL+S+WPui8knJnIuuvnWu+jDLa2elCR98QxAo959xDi3zm9uQ4Io
RSABkjq/+42rpm9MEfi3YpcLYJXpkJZyhsSWD7HQiyfYOrIWFyY9iZAQ7hiMREVM
Rlzy8vmjaK0f1VVv/CJfC7lg9QBZxoSLF5OYlHcSVZO6RbHq/bg4Xy1qnMGFOZT6
IRoI318Xl/06k1m8jPCQdHoXuXQlItDIN7dIjMGSAeHgqhN8x785wx79Cjh6SjoE
m18zfznA2JhKtvZdA5mFwu3vqMC4JJEck4Sekw2GNPUWr5GxTFmDUDvNAeSh68Dd
dF7XbYFzg9XhW3zlxk0AREMmJ6y+vYa6Odi2Y+aj+FPNWXrnRkXA54+xkEMI8eOb
5VcZ4tN2w23uUddPN+L0I3khxbPwIP3YXc2NoJk0THO2BHJ5gfecwyqj1ggKIHZk
ikxuzHUQLUa+cJpUnp5vTDNdqDIST5sEDMkr2CTskPP7IcWpeJQHubBf6MqOgjUM
CRBDHa0xbyGUDj8nCBZqjBFoOEtLeiZrKclz80UFXawWLXb9bWAwJU6hR7qa6rhf
7ih7c+p9Q2N1/0RDTcNMhSzad8A/tDtq+NS+sN1OdI5cY/T33GCgGUmB1wQLBzWU
dDPF7BB+oc6K3I68AwBT/44Yd8id/f9FyJ/sGFnyPzodqF6WHMr3Sh8Iz7BygGM/
fDc9Pqo79XwBtIZv6VNF03xdntXMEoA9pHhiH1WQJOeadW0w+wpVcmUt7La4diIR
HE4/M7fYxmIPg11vDiDoMY47YZVFNJ7nc1jiV0zZFSZSzynuTLN4yWjALgnw/yJ9
W0AqCGH31O0mTTrtV6OiCYy60n/+4Q3UzW/PUvSM2TQ7btOEj7FRgHetaV8AnNhp
V4FXGroGhzZoyMBI8ZfgqApr01aiuIx3krxyoH7gyztjM6JGaynRkvuV6U2YmTeh
oEo0eOGUebZhxM7PHqkbJ37Nn/oxEvxPH7ZwiU5cBh45aXsFDhfJMDwqj5H9kK1/
hoFF8AB5z2aoGqzzkE8K9dwWGSlJiY6QLaZK1xgC05PJop92eRPqgTkxYc2OpcAr
0K7wHX0mSDs1iked+rnTIGekKmLJkUuI4RMwmxaF4lgByUnwspPf8iBoPRYGfe0Z
k+lRK+z4I8jBr6+TUYzHJ3OCjO9HICFqcpGnrhNfBF7IPLgUarSQPdx6nHWxKEmH
Q9JX0gOzA9tQVi0k6B0GkFsoWDR7hDDTlrnQSf8SvIRf1L6knFdXO432rh1Jw+Gz
gDXp+zPhgPKN7knJlclp2B6M6YlbnnuhBPl7Y+6ZwVTrvJ9IgAysoKSmOi4hd+yX
cz12eNFJ/lBQskyQ5dJ5H5auzNptyATxCKS07HFi34LMMwla9YDebrYRx10GK+PF
b8NTrZ3UU3lOBzKWBql1sL48HA0v4amXyY5xfVNId2j/HTmGoLs+20861WATnI87
vTaOg/ZQrv+crck2ded9Z2U8zTtSkRlMiEoIDX0643+zYzvx7Bg9dhGShXm4AnMA
h3WrSdU1zAuVEn9ePi0ygOMg5DYIpk1B9k17t1rlG6Ps/gG988iWyPUfXWC0Kmfj
HdZCLeHZUeymND5EoOFnsHCr61jUwJkerCAJCB0VRO3sC9+jEC3hyURKUq15xYzY
v2miShicmFAz9XV5kjgT4zHaLBxL2fCO6brhXtJnU5X9N/8RlgUfQ9nuyz+xd047
0GpBWzkjrZHIdF4uxzzemrRX69QP65nXerxfD6cSnq4/aNweUuhSXoeSsQGx7cDv
WxNUYZDTM2Nf3GCRvOsvgmfNvPXF5j8AVuW3J/7UIFYkNvij94HbzowwAADGlrYt
hiWFgwWNofOwWNUmsVKZGODgJC7+z4Nx3uf0/qkopNEVp2hASXkox/vCyJsQCEoT
+EkQ8+jP6qPzYo+wBCVmgNLo4qXifiYa222L8jmT0kUSYB9yvUjJeQBIv9o+G4N/
7hIr6wOAG0Ope0P7jV7OFlcE9V2BRFMxR8xzV8VkXTJDEIylkWTfdWikJ96K6p2s
jrs35P9Wwbpsq2rLCdQoU5QOijqQbd5NpPG6fyxWMs4cDHYHE1qfAZ/BObBOebfy
Cr9xRwj9J3ATDKa1zfQO+eI7imtpi5db8rGh2pdZ7gYCNqq44ZgV1XGtgm7rfYWt
c5LVbki3ZWa9/ZZL8tBoVids+b2zBjyaFNW6phAJC65LWsRPmH1bbEx8jOQn1sh+
s46hJdiQUrlt3hZxy6SzajtGJtlBpE6Nh6c8T/ZW0jhXEWtf0wNmOYQPkkFPGjah
fYidciOdnVxJHW8qn+3FuV/d8O5KLGIE/BUytfxXHy0Umbz3GPZ74Z4lhItPCC9c
5UP2VfF//HG3DAkpJj/jhIEH8c4FuryN3Qi4RQXhSVE2vp7T/J0nxdET3Ze/rEOm
jx0GJpJG5cT8RPqAF76/osYXV6lZJpHbj8cEMx+UcSDMtFnVr0yVI18mdDW12ooA
/eiy6zTVK5YPpffN2H8Pmn7WqnTuo7HT3avm32CUJ0sdzm1BnPOEZs5os5bAqtfo
91oKCYY9ig2qfSK5bmZd46hig6qKH1JtQnTBb4mJpDUNX4UJqQznd9O1qn54AxhF
MHECP8rHE+SOV7ttKvAWoUvkuEx4dQi7jle1582FqA0VyG8i39t76a74VsgeYWI8
caVq7IK+IjX2kD0eIVMi5avjO8KlLxkRegAIQJQWE1+rz+nKRGFg+3YzCZS6d8nd
Le8llbiyS8FBRja2pdNX6zwLk0MHv8+m1McfnsWYc340JtXchOCSSmAJCw1GH8f4
OHYgMuXjal5SUqIm2cguo/kBCJBncM1QZJWr20iMHnmX6JZVkDjXdyArwlts94M+
UzRHDxYR+ym7L9FtG9lWbcKR6FfXZkOOlF0tDt8IVARknVa95MDVQ+0VsadepgyP
COJvI5QE+UukqARfwE25NBg8CBujPpAZmtg7R5FSaD/dRwLcXpJepbW0+aHtl6XK
MgNKEYtKM0zZI7dfSsPwijZlD0dwJwXJITz9RERlcCShUOb2JXfE/eg9Q6KjZoWC
Fpz0Krd4Owiszsc+2WJZKyV7gFCNcipbiGlQK9GnVXql99LdB3lrdwnXenlFCgeu
iFibR9j2nMtp5WZWIwd6bVFjGP4z3e4gVyzLs7jAVNQCNMmEc24IuLXm9EJ3gsC9
KLFM9UGncuYQ2coGnVWqwrfU/hr7A6AK3V/GMnW2udLykXKxAxBOQDc1w077Q7px
JzKMk0X/smtBKjXKaXT2mHjfYGuYH76HkvfSd53XunJjl6D0Ov5bsTuPWdvocCjP
KFvgqv6fz+gqkU8vsSV7N8AqI2YKUBUn6j46yG8TkhI1Z5mroUfX9cCHLyxlNKvF
vW/8a6pNE2f5BfsmYhq/a91Yud9C1c/wN1hvcI/2gsnXxgEgamjHIHnkbjj6lzMN
7o3pDSDjk/EIGUPMf5b5hDXdELzbydwhwxnDySqtJMozRNrWkBUdJZfgr04G+9MB
C59XoVqufj1VlTZtEa15V04EV3pmiuMru9DwtWiHb8amvWGvMT+ze8WXkt1y7Cd5
6cPIzpVtcRW9l9WXm4gOqqI4B3QX+lONX+2MA6lHky1LcB5v+a/t3j7HfNPFvy8V
YKtwv1vKtjlsX7ge9yOoMYeXhEtmrsSF8vtac9BVQWm01g7m3q6JtTVw8i/k6jOT
PjJzgq9mIqpsip9R0vyALGgu7Js8/eOoeerTU1lIuRbTnAHp5TSi12NE/a6QJXcg
6ZlXNnxNQ5159iHKkQzzzwFOgcUmnvZaZRQp2wA3uH7dKxSMdzS28KMg+vdkQZtD
0j/sSZ2iQvwOOTpRbTVSZF39MNfdOKPGVvCCOjR45W8v08I5vv9YQVDVl8Ki2obn
03GfN02GIHJy7auu5zjFPEm8lBVo1IhNAi5salpdmlCASJ+5fRArt9I62gr48023
ZtwBKLKzVAnUSGkBgXdvNTishmaVIp5cDa5CuTD1Y9RbwxFVhqZBWUq0g+0yYLV9
w8dnuqPXNw6fZG81i3K6vJCbdgx9Tj9acIW6ANhPmpM7AyL5llvyRi5oB4nbUuIK
VBfZTMB6mC4TUx+8cu1CbiokJAIxzv+5AxE7A5DbIhAxUrWy7kSncPsu+H7NcDNh
f5K3kJ8jdXo+pvcYugT7vK8w1a93IPNs108uNrWA1CGBjgdRxWzL84mWp6I1LN/G
Yix60NJSYxvPbP4w89opluwkUv6sfxCsYNfw+rx4UuIroJyIM4nvPN7RMoTth91b
i5RI5c0bOUGO4qWTOdg4Zupedia7M8jbzFcg41quwBdvVmy42om4LuQ6j/gX8DKa
pcCy9/hE/3CcYhUufW830QHnLpaYRA9gwxmGz/dc9otvEA25uv8K88tF9/UJRetm
bZ6g+GDTKfC46fxFjGGMnlK1Gu3tZBoZuJuZXmBqmbANP7tOTvAHun3HKFP7ynoM
vmcLHdzLuIy1ckt4hVfP4XUAmRXlNc6YJtUmLhunQ63iQ1C5F0DTf+yThMxAKQMm
ExVU0u1ZwnZ9ONAqh18TGW50hQcARNc3PWby0Pc2SvCRseWu7uQIyeq5f+DXgQFB
+FU6zOsBQ7pnZ3kF9hJaEybR6e8Fa3x98xMDPSXuBwseyYX3Xx/yS2c6uYjO/TWw
ew/zxEdCzJ+pNxQGgkR9/qFR4kmCNi75jQVcR+stX9sRdQjrDX9hmuJA0UkyG2F0
4CNm9ygW2p1P6j0dXpyFf83pPmDIckKDIUAXKmn2j4wR+v7Ix491+fVpAkdxXjez
a34syDw4+QkB2BQiXPOU60HdJAb/WAHXRWx3s+lXRm3eCmJVolab5t4lPQGxfMKX
v+HW3UWLB20EnbMhT9AYMgDLxUq6RAiZ5F06lXAQbSRri2vF19Xc8yCb04ajPEH1
f7QMtjoQzdDBTIL50JuyIPo+MzSHQLoRMe5AQVI6QfAysm33Gmu6riDBagwvQBJ7
adQmeKa+QhnNKDB3WL47DVSQBTzX/wIeTMH8qtzFxPvQvydrPFs9bLBeRzc1Uujm
viV+R/P2jX5LYVjZmTq6Bpjtg202ZHSiZhxrLh65Oe0fweIPnkHtc8VO2eCIsJz9
N6LVYlCIVvVkZc1pdfZ5SHYqfvny1aUblD2qd53abx1PjCEmnRfdc6xi/7Pjk+3J
pSDQZjIeuNopheFcxW3aBSPOeQbWGCMjaCErJ/D8EO7aoCKGpjZ8cT2J27g2uIuf
LBKeRjEo04DJKbnBqaeCjIzbbqAx4tA9Cd3Fq13XllYmWvh4uQygYIrYB3vy3QEK
Mk+1XhO0OWxbuk4lbUg5IZ8W62zC9aYKXPL5AHA76EVVjkE5ZuLSv79aHxmRFeKB
Pb2o+wXc6oWl+eolv0IfKFQFVGUvffOX5Fa591459SXRmLd9Al2UIfNi0ydLayh7
B0TEqyhw3qER7mZ+tAKboCuM0F4ClGiEeo3/OAd85vNKZ3yUgpWte1FCkSWzmFZG
KXX6LagQPwfLtPQeeqjJp81pzstCU7CdRFn5czZj0eNzgc0j7Cmjh9LZ3DVc7Kx7
I+t88kj8Ebh4h2cN90JQZbU29i/HwpbimvVQ/VjrIOteMSD+7c2g2FWRGy9yhxr0
HCoFwnIznTQtFLfN3Z5yNfpdWiWEy3LhTo86bfHQcdH9JN3dwiSH9eBKPF+9HVif
TjCKLuY+pIZpKcE6zQ4XHGQJi3xX/oRyiFwVxDWIQy0dJ2WHYpF76+T6xStU3CTK
IAWjhaBCdDwfdMfqetpvrmw/OerH/S4S2at9j0tEasdP4cVqCWTX6dCua7Uv4GkA
MSAeIpcMYo0IU/5CM8kqPBISmDp6MVv1BS8tTRlAmjdT/IwqgCnqLYpQBFkUByUs
ETk6qX/WDX3gt6TpnFFaW37ZTpmKkMF5THyRrMoD0ZSyTgFltFJz2gLffzN+59At
fzoG1/8qBuTjLF+bzdIJLp9qVR8x3QEsDmBRBK88SZgz+It5qHSqH60xFJrz89B6
3mB6qWcF2do+YLWaOITGGzkCjnJH0U9C97/aGn+FmxXLH3lnmqtWvaNgcoudsl08
VnWZhvV+eNiChr0r1jBIv8iJzSKbpTLAZrSzjyo4MU67nY9LOcMvI3aspzVsv8G7
x5SJwg/MxTnJceQskTkMKFJAaikv1pkVnPl4GDM0Kn371Z2xhCjjNz+o6JG/oEGI
OX1BRjM8+czZ8I60sNaIJnUrVEV+RK697/iF8mUUohVW4b7j/LaroX492Qv+P1pN
+SpcCO1LmRItXaeZv/mrsEXBbs6rR/pGZzx6J2skjcOptw0H7kommisK3asm9ULF
par8LRq7Un9F/MygEUAMT4zM/WYKD4rwf31Hy8ughDP6Ha5+sTDphV3u780GSt/f
O0P+dnhH99EFeuH93APtUJWeDoQLdYTuFHYRJOIegTn0SaCKguUyboQLbXCnt9IZ
3KOlpfuo/Cxei2T1Ni9hn4OYI80D2CcFp05ehZ95a6DK6VFh0+8UDZsktxiHYUSg
1VPR6OxBM90/07YgaPGUuBgxsi496NGOD/rZYRv6+VzrEQ4ADzv3bUDEHI6mjxQ3
vMPEj3ytfMEDy/WOWUO+WGDGRphBCnjlb70peRCFay6mFrbwYP1erXjtP7T7bHWh
yKUUSW/oH5uqfIgOou9/MuKBUgWhVs6qTWsQZKMZl4BCuaVeJ3rQ/p1u0fl4Xojs
9JV2Uy2XlskrQ50KBzE8QMQ6O04swtt0bhJ7UzF04hRZxb8diGT74X9MlaQ0IeKy
iq9Q7PEADS0pjIQOzmpQHSg5gF9vaQwBafabD79zRRadlWV9jKykHuQazFuQhMbG
TPVhDaBapKa9JaHmGRM0Z2DRTPEapcN1f4487KBpI3BSpN4TjBg4b6FLfVn3p1qV
4u5MKwhp/0Xp9RzeU9d9eYjgxaJAqqJcZLQqlDDtas3BWzx2RkCTxkXDlLJdvkwS
bt772vdHlkg9vDorEOaNlGLpM5fm8DR2pe44pqktbJGN5Y6MH8wJUGpwz4yO8Eo8
fFhRZjr1XTAL+ILz3qbFBGEXHVBCcsfaK5+luw0KeZx+R/US7DzMnJB8EED3f9lh
LR92jvRuZ19gIpB2UOcW4DBuU87PT92e286Fgn92bNHH2ds55vYDvCwH0Bn8jy9L
wQST5dM36it3LFIt54biTdD3vJfdUcf4kRxGXx/KiqQHiaAAqY99a+2uof1C150f
FPr44aygqzVBV0Bis+6jYaS2oUZQGQOs10HoClvmtdyrSSbiRbkoTs/lIL8Ly8Lz
9qBzAzWC7QmhNbNK1iWKOvco3Ck/LAuEH+SNHpBXiitEZ4pjjjBbUb9ziOaBaVVE
IKTA9H5tvENgGn919wiv/54ZmS2VWTy2+gPZSr1mPZAdrbzRK2ODT9DitNhxQX+C
Bh/O9O8m3MVESktGfiziv9pNfYOcRladfArIUM2YsYg639WAjJnwX4SxUUnX7R6s
Loua/FiiAd9JcUMBgeG2fjqqssVF3VuOtI9/tsnzL8Czzpu5A8G3jgasNY+VcxNk
hLEulAS0Io56i9WhslrJetFri1aPfxo98il8h/7mIHi/pzfJKpnPFbQEeQxcskQV
KdSzLlLZ1/5PHJ2t0TN3m6gT+eun3jrW1RTbuv+4RDZ3DHcrR288g75s10KbgnCI
NlmLkceCjLZxtPUKyY0sBRFz/3VPM9QKrY/9CFusI9PztF139xiWRAQi5A9BsmYR
1pmyyE1fbCutQxKpphLx+kzpEn1mVK5SmkuT4YkLAsJVrtHQh3ObeCJQWimymrR3
qby/X07zq4gNcAtb8pDpDX6MgRX58Seuq3kfwDZayILy5H/Bp7yHUJGi8+TqDS3N
aXq3MHpmRMaucByI5JfhBPENl/NTeg9q7dURHz57iM1jLSWEuTwbQ1n0QzvFKuBr
7bZWRXEuua1GBN4V5veWmLNajfJdBK2wsbQnDJKJ/JAFiRlbj3xBvBFKVpwjKjGS
HcC8OGmHX3uVmqxI8tTRFBpdk1tl9EMusCFT8sFJ4mBAwxgSQRj8FCazyD/cFSmW
ESTowIyc8rdFkNoM1g43PcSMsEo5UpLlnDn+ydeETuyYJg7oybb6BMnSq1uLcysn
o2b8e0dJ6Z3VOpfD5wqsV6IcGoWP9Iob5vTzwqZaTaqfhpCWneHDRKlxdaqzyUKH
JkXnZxu2EKkzujtAKH5PZYCCxGAgcPF3TwvWvdtGrme/mAfuVxxaKapmVtrUKPm0
140URS6p359zjamaG10V+vnHIYAHqDl8y7UJq5f8jP3gP69VIJTsP4UMsZB2UsWn
9Pxm/iQjpqFYjkazP9z9aESKQ5KPOiM0InhW6W2QMU5bKiRFDyQ53+SqcRh8fQBM
tTfnz0gY/u4z2RL62SHxRFcFZgTEVwl3kZ+csb84jzCv2Hq78jb7URU8DXysEHty
pnRLD1wMVqlEGEZ10ddUtlAgMOh4ZA1++fRXgnyp0pAhfIRi6tSNAq6w2WiIc8ir
3xm4djcGSVEBlK3rLUYgo02xVulOOAsJgk0eUPshrBr58KqKeqgf5C6vDp+35Nf/
39FG3kDDnnLtZy7aG9AIj0MHMf7oX0oQ0HyW69Bfp53JzJp4XjTJFat/si6NDWkf
xmUeK2o3HKGkXF9YJdB03ka//5HJxQAvXc1P2h7nVSdT1p9ADKST9AjXckEgzBU9
i5ILLFuZWCkM3Bk6spHWYVChO0WhtuyFH+1KeqBtg+BY7lR+j1Rzow506/eIOdLz
8ne+8qflMdbIMzgfxY9QmGCffUhIH8v22/bCb0DNeCn7dIvjmBJPwbua6778brjk
rtKk6jox4ZzuKQfri5j+dbvR/nEu+PCHElqQtPlS4+/7D4fqtaF4O6L2LZzUZQpE
tTwO87Aae2+v5o79Ot/yaOHpB7jkwrCyUXgByUjQeTQ77x73kMtjmk4y/kLPHqFu
i7RUvs/lF4SVOdf90dT1/dqdUtJz/3BKp3LBODbwBL1i3DNHcCT3r0h2vapyChRR
lmWXrNMZa3y/O8GC2MBzGMUkLjFeicA+dF4IY4thrn/LHcLcr4IJ2bJttYZR5+Ak
R6aWS1q3u9hkwShjZ9hjcodssd3oWVxDanJFxbSNQFmG0g6sSgHKyE6z2gZbUFYU
ehPUJksCPdi0vLkfcRlVQo/SlLIHSmFp/nXJRMHSeMRqcHTyc+/OaDgx/vgQEoYZ
7hEwxFQXtogYoV95ZWtGWXTZ63WoOZyJ/Lwflu4445A2zXDZm+o4jBAOnsgst248
KPEcBzvgH3HRzhalO96EoBpxDr+Hrkm0HU04d9uEKppwJ0EZnQVa2WfpynNX6ryT
PJu6YrjoSLvY9yxohRji0ZZESortg0tBpJIBzeqPno7+XwrKHNpQrZT/JwRjbZoZ
dZc6p4jneKC0tQfFQzsRoVjCZN/OoNZT4vGNWgsfHcuSO5ltlnpJfLCKQZEa20YA
4RoYIrvcbcr6qHGjcBD122ttc1mzgJxdpAytqBmxwaHmJiXL1KHHnPQXOjNiku9k
VunAVR6hOV8gxQe4QPgBwYtKrCjBJ4GE0XKi8jLWWeq3OtAreVtT6WQf7b1MKNG1
9KaMEOmjhQioiuyjdj2co6wRUR0UJDV5iFptRJUvwWc2+d+XrW6sue0HxTCF9yMR
ysAkfTP3AsjYlATLLniCHooGYJkk4bjURY3zIcwO+vgoOiPy5uMt33HG6Xw95KEG
y7Pl7eUbfkMg8gsg6MaZXR+N70w4zEob1oEBNaMofUGgj6BPK36yw2AhSvz3LQ2M
Y4rSoE1QD3+rjpERTh+ljbV5tYj80Hqj3Toe1V3oOrL5SrgXrAV10ld6oVkRM1sN
raSCO9dSwhawZdgyPfHwHBIt98BnFdc9RarrPfG7c/ZwJzZP2xHmsqMvEF9MIe0R
qb9dRYd2Kz6yKKc/knjjVoeo0oSR7RovqnjU6L1jsmWH+pPXbzLj+GxTnfqR/Q7n
DyYWowKLd3FlVyJXCF5d+uV0F6QH63mlduIDvVb6lXOlfF7+fmnBbUKfEKefdyG0
sSaq9petbyAJXCikXqsTswTpavsh9LF/rnUzeCDsGRHtsaZSFKMSjIifn2A/j+qf
37i3/Luyj7IMDkK8ciTbpkWgq9ramcHvGCU+7uTEacFmwEIOfrytxqBgvEUfrmTp
iUcf6oBC9yl2tXhPWGD7lqHsZ6IJX9wI2G6mpXYTaor9VGF6PucCvllfq3aLAfD4
u/O3g00LraejbCAf6jwBorKPPuzAN7gBTWDcFHQ4fc+qIHEWIPyNLnW/24plfiOU
dS55cl7+qfLTwCkEuVIQNmWW/EMmfT2lHJg8h2hqBdVU60OV5+Gdu8Yl2Y4fFHfN
vCfzZ5BEsoJvzMvAOyf7CUtKF7hiaseHiyCC31R7gOQ3vm4Ud0lmy6atrgCvgfR0
9iXCLMBn/GNLn+6A+vaZY8mFxG3idkka1cDLSS18K9sTrHGNOpHVVoosP3iKEgaW
9O+ezLxbpJum1w96PHIRtLRMgStTU+r9wTfApE2OusShW/yDl8eahCW7tNtpc/4w
EuljWFh30KdOQeexHGTGa6i0c2anAMeRZAv/67WOoeInV0YTbHfvK8klFr4E6EaN
/nhextgTdZQPmYrk1m0Z4aiTPq7FEh3vU4i6lvF+ecoYtoeTjV0WumCYUCGQmErU
omVIwVW6F6lQyhbrMaDHPUh5I34qjbiaruP69JMWathrj6o8eqiQu2y9XNrhgASS
xKi29lQJMDoA5y9XYvbE1JJdylsu6ogGucf4xqYy652aHBZNcn+PQxOa27FjP4T7
bNMo5wdKbKgM61CkxclU1gwQgpFEpevllU8lhe1Gelw4ZEfHnfv4CoVaCv9OMvxO
tlN+N5Wc+0O8udtJyqaSGXnQaMRrawuRs6CZOAQnBqhfJPLORpPSVv4aJ6YJlFkz
FLkgubNrZ/cFIEPTvhGsUuWJProxGzf9t3d3pVg5P4jrwGK22RxosM5ONwNqawSf
enIZPieV+GgPsPKETYHmlnTlH0rYhwXfe6NSthvwc9pQM2llJBRvGoZ2ihUmCYQe
jmlBL1V4dAQrV++I9JX0UUK6UJ57BTvp0QzGBwP4J0tDxgHfD7n3hao2m2+ROoFD
mCh3i69fCcNdlxw7TeuBOprKnyi7p/e7ukD4xQZb9GMeAv6uvaVrCEho9Jsf7+yU
N2YaTiqBrYkRbo/Y/ilPYOlpreGromWjPwpzAJ8t0AyLCFEy+hPaSmCdUqvigqsP
ZlWCW6QJ5P3omAXepF97NJ/1azFjOCVVy2xb9vxzLkDb/UZRhUk+m3GNumYuLNnr
FJz7b7DOqIE+q86yVEfyMVPGPX9TeC6SO0Ys2pyLbh6CN6pHNnYSOBOWyqQrKw3x
nGcv+lOqRe7o6w6HTQpbQYbWInvJv6g3Tsch1mi/yNUWZ/m9oAQp+1qAC76aSVGu
anCmuv9c4SW6Ik9raWgvKjNSIQsiZEUAsnOKGiTaj+0hJjUl3rRhasFdM7/5/X9g
6wltvoz3IK8d3AzhgLF6Za56bAIHcic4WkTOYQTt8DlDyANJl999W/kqPlqac9I3
mv4v+amas6/XI4dWuacUaFkwaIfPlXwvr9DZNhdL7ba9oJxtsmoZ2/j1kzxjJ0uN
G2MWRXGnndcKh+zlHMwal0sa8qPTbkFIbKURo5gGJ8SVwc5DnyX9pd6bgckBLw5D
8OO4tSyYL7nRDP3iLE6HxuN3+J5wsWz+FfI+UWeNT0DyTYLNn9tIhSWikbIKMLlW
Wk935idD1GGX/xCthMoAohTIi1e+GbXt8XxR77bTf5GK9hVYAEXPovDVHL72rlUM
SOF51C8kNpsC+b8/OcyKLulWEokk7rLsd8AwGSE3bF9kfZFae1Qxlx3+swFrR6Y8
10EI+b5yTy3MrrnZgTVNjOkFL3cTqa+wr0phHUN3PNst6j7ecfgtGng3otHGeyPT
qJ1lSUclDOsn/f7iX+GFaQ2tuAEWJTonz7aCrcO/rs+FR1R5v/KXaDxelK118dRX
qFWNEscbI/MNFItIC+JOunbXU7YE+X11GY2mSAfcaQXc1KgcrcJ4saZPDvDYkJzq
jU395O/vgFZ/8sjqB20vbZcGwwdEgseWg950VviHkI/gTJdIdCI1pWitXnh/QCJZ
XBvL/pYIsrhtiekzn9+Hw9eHtfxKcBQzcV1NfcPrPNQsMkwz7eCq7iwHGedsPt5T
SyxnuRiKgyEg9RBCi7btLjMAYnoIdz3uAF+twcXMEaib6xpI1LBZq/fCfJFjRPjU
MGHyN+Gb0fXoxDTsMQ+4QG46y0te/RMn6LYB/XIr9vLUn9jcJSy7WdNURnh32s2r
aJjY0HAlJ7H9sVGyn0qUspMMncoCj05/eAZ45ycA3JcvluCAlcsn9OCJFpvdN/uh
KM03nlklBGnWc+GdfU9hkOQ2lO1A7J3mpHTmoBg6mdZh2kARou9OVKdVbHtQ60VV
ryJURYJGoVjW56JZ7qPwYE0l/kvwbH8uTzLxRxaMg8HmUBQOag4bPq1MBlXUwhFx
ZQDo/sRPPC59m+GihcASfjFGwW6oAg1ga+IW/Nm7tfsPszI0Upfxi7TtAY3TsV6w
zN6o6YfXBZMr1Chq1dzLJEclybBSTGqLArXV+8QApo6RzpUb0G0u4HhBEaYuE44C
Dvxvwd77dKA6hyzNgD1ESG00GbD4CWRDxABGg5WJdtG+ZROfhuj5cEOuQ7w4d/lb
jkjmpXz0Mshzubb+jTKRWrTwE8b8jCI3DkfBeQjqIOXMRUy2lUlGNQDEI2gzVkMo
Vmmo9zNMKuqRMPUZ4YpL3F5hWW12Jy/PFN9y3olQD3WygIKiAENRxi7nGNXYro/Z
Nlqh68jVJ8oasw94cgWGumEdc1X6bfZV97KWt2imW43zQmM7EnTx2S+0GF32Ospo
Q2PixNxEjHbm/GT0Ey9cW4nYvFEO6OajXidhY7V9+cPjIlY6N8wXHzL26zIT3gok
a76jMK1Kbbh0dtgqZqGDKOaHLts1cm0vbu8bR0SxeTJ7WWCp+C5fJs0tF/F99fze
OGJpq2RtWwFHIFsJfDF+0SKYCXbth/06gXB6MoVG2+jfmlrSwqC4yADgIyX1BHsi
yOsxovA9k6iqi2NZhC5m2Ay69FX15w4fslOo4bky2XebC/Hq4N3xAGIHSD4NDrQ3
6JNVYiAgnsmTwfhLA5ljG5PT2dZCcPJLiqbRtmn0J2ryInGFZ5EvW5XeX/jUvSwT
cWnHlUTn4bKAX6SrXb6xyHmLqDzoZ+rkRF/C5dtmXf4to77K1EtLZlP+cGqfrW7c
bmj5focFPPfroxS+pP85SyARup+VV8vKC7+icLPPeKUssG1Bmbf1xkiOVWmzVU7u
SedVbBg/9ldIfZRCeAttuh49vHDVJNG8BCcwWMsTsEJ7pXJ2fer1MQKXo6qPRXJ1
i4Gq3TlpXnQ4EPDnzi2EmAwHA6VLg3t1ruqRW/azbTBxBvtuWMl2DcyqEBwvutnQ
KxB0zHHkLeWWPc/HA8IhmDC1MY03n7gqf56XrSQhJtzwXwlWVEOEuWH0bgT4Sa43
6SRF4+K4p8pwQZefvT+TDhO8lruUosUJdi3QwzA+AxVCHwQeq0T05hgwxy7xeUAi
59eR47AWs7mKM+wYg74p/9N4s1tQjerVRIhI5Rf2ihM3Tg06ItFd3yjdM+Xn3ahu
IZsN5nPNN3SbzgIcM7yM6ll7pS2bF5RPtHIT7b2CV48u2IDeDgT65CbgUZoetI/k
XxTJa6zqUQPw3no3ynA8+e9VPLxfSezZ/sYZD1U45NIImOdrLuZAjOMW1mSIeNQf
B5/3dqxpIs6flYNVkYnZZbLplC/qNYGWZZM78JkNVnNYVstccJA5pbVeNA8ZMEoM
DgFq2dtbqExxxwRm9E/XOYcAMTHFAJCm87CNi06Pz7+7IfIKvohjj8uN5dqOSLX1
kMJHnsze7++GqigU8zXrfUSf+ATMOHWJ5JDkeXgIEUroqlsp9Y6JsWRxrYdaI88Y
s3T6SizuwvEDMQ8wpN+uJvNvHgYn/YFwH2fSF+ve5G79XtFsqQq8Xtp1LflhQcSD
XmI5RWWqchIjutLa/vRB85FDECaMmDqdsKFz6KhmQlJz65zmHoOi0C4tPf2d8ydp
cU1ThYub8JsrfgLBZSeYT7CQLW/c7hg20XDmpPuLpSS/4pVYN649FbpiXKmEcaPy
Gkwr8o8zdbo80EAUJJVWBsE6DNSUCkYl4CK6VbviMZ8hLfs4CN6J/IRPHlqLDZEm
gae8oLzBhSdf4ELMXgCr+lADxm1DJNDkJjDfaLUmMDobKCCnwlSLOdfC+8E43WFt
fbJetenN3+ZQqvI3nHL6m9jGuZ8lPXqd6OOGP6vm5T7pldxRlGNj2Qg8Ef+JlA4E
nSwUqsGEV1wIipcWBMSSNot6cXiBOU4ur3GLXYUAAew3J/Ihba/pzMaNeu7e/uRl
fkpAIGWHiypC5Kb5pOR9arkkYlGAELjeMSZEgjakyyrNJm3idqwxZ2bOUQVzz7MY
3IzOvOoseuTUnl1DTUncaaNbqGwgJ6enE7gKBQ5pvOdrXBl58rcKFXdGM0prmrp1
V3T8B3H9YoDJLLZ6n+kdk9q23DtKgP6D4HvwqcjjqUg8xT7+kWz1MgevaMjeEtxK
lTX9NYXU362f7B2Ba4+6A+OG+siUIvCkCHVd1teJbtvMFNfCSkTQbaq5mi/FG5eQ
24DNorzVXdRC3Iwi8m0F2fiy2Ku9PelUkR+T79FqX9UQWppBf6GxBVTe4oV9+8AW
iRrQARt1vykdhuwu5c7O2fiUAyWYdaQ9uTLixT+VFwZfnNLwmQdWTdHQ/YpjWH7x
VabLvIHa8mskqjc5H08XXsKSFI/MfK31aSxy2HanJ6yvM2oQM6ocZw/MdHLMMt74
84O/pjOlzJGW9/3/W8iIUe1bZuekDoywAPyD4KaNovEGnivT27qR1OlQfoqcEhre
bplDT6bSHnanktUU2q+JHG8XVrWqpfvAjUYTh91liRFDGyrw3e0o3CWFi5/9GJ8t
4rrg0O+rbBxFfAb7RpRWEgsMTp9upnTqnY2boYFSIcX35p3vuCYo8Qjj2DgSSBJF
xDGyeYj6kWTGt5eLBxOrLid21JDqpuw5T4eXaaVkykdd7n+nIjYc9B4Fpt8L563Z
1eGBrfft7xVeKbgja5mObyq8p/nKMIshscDvRALvnWZXaV5SQ5kHe1AM1KhW00RP
pVJqqZGPAd2m/OfI8lL9+M+N9V3SgvyUxEtTH1H6GsDrqH+btM/5LnywZJaDLw46
z/vUqMZi+aP5NZNwdURNRuaQXZX0SGe2mFpYopYYP2LKVNRNC6CUNsMwbvBr8B21
1xSDPqtc4yvR0LHBwRp/IvuTpDYVhXhVcF5639AymJmaOlf5DjlVptcr8jFu+g5I
33x5kz/BPeIz4A/GI7xUkUk4X7Qg4i6S1+QS31BWULPrZVqgUD6oI7FWY+2RQhz/
bUmFR3MFyWT5k7j1XtF3Bl3prNhFhrS+SeWUSj7AELTYln70c+v6jxb3MdE/oIjd
KoPc7bzL8Oxcj6cSV007XF3K/qReU9c+hQK+jamNSp9QXzvTWsCwhdWGy5IyleDr
6A2wy5AegQoxuHO/nKxq4Bt5l5w7GG7oKje93FXiElVG2l2w65NMLUNmd3kAkDWB
ICyvxwv3teSbRuYogvYRZWPjhR9iVNuqYG/eWynbalRaFy/G9Ewq/OreQbImwLXM
XGZhczZYgJq9leuA0HlCCtCTpvaFJ6/RYobBa/ufkFNYXqVkMHZSdsaY/3IU6oUX
XuKc9s2J2VGJDB/ceI+N1PILVMgcubNP3CyDxhHQ55iv23Q8aWbJCo/2CvcFt2mj
p1Z/6yw3Xvz6Zvw5Hfhk4RfpAz9u5l97F3LEGyKDclNJLvRxntH7w4V6Tlp8+Xno
aPg3uP8rVoFP3p2GEoK/0vgY42T/dOwBGiIjodXx/pPNIuOfxdBXElv7fXhYpkMr
sm1efZ+G2h7Kpz93Zo0es+czUi9JjDscEzlGUwNPfBS91y40HUR6felRNJ6eTBur
wlQa/nRjuSwV6rjb5rtNPYifD1HNglVE/TbYHzD/n2QE2e7UF8R9igsg6O1x+nqT
gwMBK+k5oBHZIUCF9b/tcx7p8CG7fQvycQUGmQe8PrEd+LE2iVZc0ylKaDp3+Z1K
JgcEmlz95epa3ysJ6diKBC2pOU+ndSiDzg3rH3aQ1Vs8rIosvux5GfFsbePh/Lmd
SAGE9lmGANZAen77GiIrma5OGd1/ZFTfIOl1izLruyx9XHjU3RJQpzJlj2jMy+nK
OtGdNwNGlLoCCePRGXfhaa3upgbXgRtHA7vWMXwJfHvlSUCvDAFxmpt0dWvNZg7h
Pp/MRtqRnHKn/Rmvz5NDzzjsDML2ib6yOSdgP4xQaZrgCSxxCq46DnhicC74tMc4
/ctJJPUmpiGR3U8MXRZ35Qg0MXdwfNp8ntnmwNwWjLHJBMAV2RA94uDhBZyh+W4Y
qF2FH/0mqyxTmnA27csB6Dj2B4thoucVKPJPdvDOJzZy231P3rSE/EBNTu+7pJMf
ym9j79sxp10sm/QjwMUVOhIKCw811CIHpw4/OBrnn2YWOnoAQf2tWRPfcemAN+3V
SFQ7acyVMv8ruPQR1+SAKsvzNGhBBh0uLydnusKvh5NANX5yPpnYlpvhbk1wnF5p
FK89IuQt+eq7/S9VCR9PSbRXwVSTveMFgxqglpaoeaFotV20rp+3wBTbjzVfNCi/
Ge8onMrimlaWjShA2oqlolNztbLptuRlOXB0+YB2E1uqqkdqN47FE94cXKDX/YFC
DDagOxLlWRvaibQ4hwVotDVqMI+CjbRu1Oyi84i8RWRr1Ub3ckjZQltKoYrRAis6
TlybrKqzHEK1srtO5BJicu/0i4RMm8wFGqqbhlcVgSP12kFy5k49z1fQgm2/+sGE
G9wS0mKtnemkghav1pwFBYLSwHapLl3aMIqVLEJoIznoO38aS044p1TAkTd1g8qp
+f7hjQ93/XnpAzm7EpCWKn9B992n2ladfA9IseMD2j8b/eb89Mo0+Umqdl+8bZRa
nzVOmrXaPax14Ws/6JHoiY4od1TlwaAqoWX4Ir217ZGEsX6QM5h9f/vPEdQre7t9
dcxg8nfVBYUNZGrY1jkJDUrNPdsu0d0vXgzb00p4SGAq09Lof8DPPX8cX+CVP0pi
5Q3PjI90R3oMhH4X68A4uqYL5PCShxg2dXP0AQST8lHTTWw+TgD1IyztaVEqmr+L
tRH1tCJOv4hnt7q/X/ueWLiSyqSef/kTmbsZyvk9jFUAY0jcHuXodi9dGTmmROc6
n2y9dteHg7sf+XoO+xYaMLbATfRjTaYUYW23BfU0hAuV7IHS5JMTuucI3/7Mg2ih
wXCz0j+noHN4DCrBW4HDydprEycPl/+qWCJ8zqwKWfA/6usQMG4gv5xjsmDJZPvq
gblZrH9o5O2k4+9S1VC/nZ3uJDDjv4tiyJc4EhuEQjEp7YUVwImeSETWaB5O4KKm
vdOUY/NX7t398PrcXdw6e67aJ0KeG1XkpOF3RxNuL4Oj/nsmICowPfcSPRLfOYpj
kNz/5+voXlo43Ohd0eULa+JfoBrkK/osTcZkQeXnHPKKjh7VbdOTnkL5Qqsqw7gU
V/7NQeci8bubsM5KD4WCca6hFRgbtY9atQlFG2D9B8fHp6lfKdBwENqsWEY5CwtY
5AKb6KmbnchBye+VU1IBvbq+9+2WzGisnsI4T1UpP/6BWrohu/QDDda2IiBYxEyX
zk2Vl7kU3ocNiJW7uvweMwdSPH+JD8EWeafkc93HhA48iaZanX0lW7sPuwU8vfE+
lEFE9hjTeA7TwXfVNvr3YtqAwYF/J8B2xPA9RTagVTmQdb4o0exFjx94cuQ8NNVQ
u2a02GigGgOQvTSyd8heH2jttU1nTZJDcWXZN7i9SFbMxi/e27Hh/7a7e14oL3/2
mtiyaZ7oR8UpFZwPzQABVtogJoyYhuri1jMqHFT/q4SK/ngvFp9SJpuTBB/OzUyQ
2kehLr0bxdJcxmr4vCRffzaZMKuDn+iM/ZvSazgtqlv0nWs4Vm0b1evgiNFaL88S
uvfwQX6LIgtKrtilHlf2egUDSlg0SYGuXRaL2aFRr8S127n7IekM+mfJW5Vnn6sK
wBVerd0JO2YjHVUfDdaobkU30jtBFrc99r1HzKbavGdM0iU8+PJk1Tbut74CLsI4
TFZC/gfKp+DOsR9Az/I1AZtPlg1gYZcY45Sy6yPGX7q6J2W623nMv/2Lex/SOfoe
yiVTUsz3B+hGJQDp/zKiWOyqN0kOewt22hPiqXwHbxAGgmSAR2dJww5v6zm/fTIM
2OAu+ikspIGC0KrGWCq0OhIKWnyWBpsKBwCgKumY73pMC5fllgQQZX9GQApF61qI
rXG7VfMj7VwEHQq/Z9BkEKvKTMbNFCZtpVTgbd/7xBSd1hx90g5Fl373b3IL8Bcu
lKA8PVmW6gVnMpl1ScqHHR+Jnzk9vPVbtgxZ5AFL74cs2X9WRfftHZF+L+2njLHt
8lsxeDTwmOZ1i1rPZ6wkCa3fj3jnX2ps5Q0BTg0stz97Up9k+kDVjkCur6UEEaqO
2wJjzTxBqcQN5uXFTF338bFtc8Z5XxWoA/DST/5jtDg/VcG3l8cAgBQm3lZ9+O/f
cPr7go5hrr/ZdiLPwY7YTj/Qm5xD/FsUpI2zJIlFvSvgP6z8HEdyiIcmRcBIu8LI
z2ARPy5iZfJO4nQjhp1BWUXMA7ze6jv6hKeDO4lnhP0QwysOCwqVC4xGH2UgOtMi
kzrZBA6uSuQmkrIkEDCTh4BCOTbvYCz707bZqZZSnmZQ2yTnlLmZonhmlgJ3BEqV
WnsBx5PQqXQ8rpAa1qSUwzcJ8Jt4YD74LAPTL2FsQeCx+rlowBlx2F2+zhM4IPR7
QmL+hJIcNG0T5XGIV6HeHE0xTyycFkYkoZqlJCfzgI8y//AOJX5YKTQzOLKC4wnm
6cWGbc1O/4S2A57eiPtokl0r8SElLb9yphg7fMvOvUHgVkibcXxWZDSaWFNCSnZa
79rXAZcTo26BDDAsviUy00823lfsY8U+XDI4jjJvueR3PHiWFz+Qm+e0yBjJtFbw
BpuAzA1OIrMh1j/cVVgyN+onldLhEpmcPydHQoM9z7Le4PLBcx43QfNxmKASrmOl
6vhcRSfniW6R+/lUVqBcM1qa7M8TvOYo2/0nBYclohtaYw1q+x91SFOYBlgyMJ9k
Yw/kjdwJWV5CnwXhqvddkXkcJo9JqQyBitMMramrNuw48qVEaQc5oViLKm8xgP4e
WG02CmjlQho3eU3IzoV21HHA53Kb/kA50HyNj/Lq6QkcWmwuArqz270Y3Scea++J
PqdeVdWx3kNxCtslUT2HQ4Ux4kdEIPoBlQ87lyCojLX+DUJZUmGUHC4KXGJ7o3S5
eZA6kI9n/zOtpsj98LcUAA3wLZwvtfY924KzbBKuDke3AG6Yp7N02Rdd+zKcJ/z5
BVsa7eTwUsm/4nVfgP9qBmZIzNvyxeJl6qRhC3uBzF3UEaIqxrQ+eUUsafIZdbxq
5LCA3H9dtR7vc5gGFZCjp5uDGUsrqSgZUYmvrla+2U/cbyZWDyTNHur5Q+ExqByw
QKjbzNui9eFyNg+aNKG4Za8zruqgFAVG/KkQXdE11UqWjOXtmvuedJhcSnJdnvuD
D7BqIYdLD0rprrqcQPoVhTDFchmaNVnQNpXB0Z3qk+khspw0GEgz82l0onUBwy2e
nvGc+GCWlmOVGc6qEV5Leunv64y8faUo+o4InCCK9lRgPsP9xHwue9tBZA8Zhl8S
7zYJiKZHITeFCTmxmFWBIlmffFeWe7M5Jb1ju17DwzHp0sYhRXCKMK5Vq1vgo+De
JMa2LTSJAL6VeZ033g6LEI4utikU6HrN/7Bz/6Sju3YfMJFnEM87s7O2fAqCxIGl
RBKi7scMY/9IVxVWnpuwycireOh1/k3UCKqgZaOev2YzVjqg/gApX6kbAOGkS7Wa
DlHwQ1cVE/X491lxZr4F5UYtWa62kzeahL9of6hSr0YILMhnHpBYYLk/WKwRhfB/
J0b1LapPSRum6v103h9zrkdD4bp10RvX/SwZ6BA4XwLg/0B03lhdURgirDSquy/c
/abhB5MVh+8mf6kUQPnoDwc7qas6nyfY7ZwUMtyEk4e6zUp/yneRWxdjuZSPH4hl
BNVHX/INijtMznF2l6LAoyQNtn9z6o6hk5Adg6cmeEkraK3sji0qU0DRMLMASned
XFxoVOmiWQ7H5D7pEIRW326LnF5d+mYp1XNqngQZKaJ2K00KmHDXHInFvk9RLz2Z
XSsYySYhFHF4V8rbrdYKzjM3vPcdYTWmNdQEX4K8eOUPZRdZFeG3/rbDnU/9yPbI
uKj+yg+AuZb96yGyWZuBCVo+tLH2XOtrk+VM1wGCX9JjbXJlP4AOFKqz2+vXrD+0
iWCg+2p+m0OCvDTN/AqsbK/kMCMJdpGEJZLjIJbB5x/TTLl4/x8x0odjeKrjokdM
Fh4VDRX/4nI0mZ2G/0ZxoqxMUy1KpvDCZP3F46+4CgR0f6srWAgke4LQIpuXas2b
we7EsHfQDKQG7D6k/Fna8YEgqHQqJuwS5SWzShreVtsqVrrU/IdW76Cv0iMW39K9
6KrWiUD9o+IBbWpFrMPBamLl2BuRf9d+UhJvx0i/l3g9T4fkffvbEWblOKbv+Y9B
15BFBzohDnJJ7HlyaLkqTymBkkg62rE05Y26RLauYsI8NFHKAPNb/xXSNklOJSJo
vO+s1WryfaBDgkdLWrjZ0Vf47s5x/eYbr/5DX4CX/ugJ03814u3pyYb6zOFKBDCn
JZD0y/ffaeAvVnmYJVDuedQicjt3fI4l1EYwhC8FGjFieL9fCi4+3u9m3JRF+0kQ
bbohPXctPV6kefqVGgC3g7oYKytKs5cci6fqr3uNHAmtFKkO8OmurfYNEVKgGO0h
kut2+dGz8mTvHHGwMONh00xCLBo15MvNfHCIHNojSOu6EyFUrmq40dJGNEBvlyUp
bHf49XXn5JRTl9lhcYLUHtiQfBOL5wDhuQ559BIWRZr61NpCTw1dfl8AGDc46qKX
OtWo7Enh6AuvO47oSmZHa1cQPjF2EeLkOG8KfYp3l3eKd58OLL1FpjXxsbt8NxAP
+QMq8DKbBXg3Cx+wzcq9BjT27C6u2Xz8lMkjkVjOLWcMByD41j3r3nHThZPQMBPM
9rEwktqFyXdatFqxAOJU598xDcgOukns8Q2jDPxEDx+XDLjEmziwkbv1qx7ivgCD
lEjX5yNpWHpGJDYxciAMIDkDh6j+/swVtfrpLKqwnZW2oNNP/DD970HmBhLLcltx
+pmTK0Wr5f97b+AYE3PcJMCvw6/5ULEZgeeRd3eNbtoAMBTOh39rLPEDPVVkwrBe
lgCbUfmw1ljwELN38Dp2y8J333gQfDT3aMSrI6mbadKbGF+s2Qol+nyaOkNVLEJZ
X+gSb1BHDeCyfxO86fHyMZrrvBzXCHJXnYucChQfd1XLEpi9Q/pwexyXeTe5R7H9
ba3cPrnmtZUj5ywSuhYWB879TOddx81eaTOHZ8ASMYAkv2QD9r+Vko2ZGbuSM2qz
cRS9llD7LyIfn/uZGtfmkVeeJRqeo4CrVU4/r+Eg8DiCeM+ypE7qwP+YWGL0bUR5
Oma8IWMZL/XWiD3x7HbMDWpb9YTZYLmF/cdbr4JfU2o2k/KYAU1k7cjXnxQNWIlT
7GFv1b47cQuMvfFkYyVo+ozGtJGxrEwQG81TPChC/ZMjnjogZnhE5nofk4nkR/UD
LybKygsszbRoqapN7NbgJCDp7h6/nfk1RSvcOVFN5NzIkBxVB8qfcOofgp5Wb8sb
xZtw1Yk1m5oCoS+St3tEkcBEdK+44guxYDZS1ghcjyJdyMzMLBfPv368trC6l+85
J8y9kAK8TUS3Wr+tXPXRevUHXtnSx5w3AzLgdSIrrco3lgXAI+qb9337gyJ0Q8Pa
KWm/+u3NPON39QSyXgZ2zz+35PCbq9RjEXs24lrrsj2skL47/W9QEFdSpFALobAW
KmSWC63XnzbZDf5ww9IeQnsI1VwwfJhboZ9PGI2Ory1z48V5M1SzkviDZSsFBxCF
/weteq/7EcSbESXghLLbFRqpJgscAtPkVux5O4hbxURVeX5Q5Hn3QG7GER4ErE95
rcAEr3xFUlXjQp4G9t2bWTrk1OZVVPmDp84Md6d++L9kJhXZsQsscFEB6Go2iNs7
KKTCYQ6EQIvrySw43LBeW1LWNs0eDs6wq91Dsryjip7TNRjk4yRBhM0WMDILYa5r
P6f0Q5frh9Pp2xCJlQLhFh6ibEa4IOacv/tEBxxrP99r1owkCZR7Rk/Tg8pD09Yd
2nR/u/4rfWUL3VzFOaiCb9HWKiIASaNDOOii/hpxnlHTMOoDdvk3VKemYdx8z14H
4/0OJVX481zicbFna1voTH51UmtGeSMwLCozX6PAB7S1WwKNVuLobG9y+YyDVSsp
FckzzUaI1lZcIMrpZBOp3Cz1yjyrit96YMuSPDWa2rnhsq0BlFCiCNHT7b48elA6
U4hEoeG14okLFqXH5vQ0Wm4PgvvxlSls6rYwOVkVsC8rZhG86LgHb2hDiOQ9UZv4
2BzQJi/F89+Yy9W/KrwKdunR0aS/Bxvk2UnZBDKhS5ItzUzOoKNjC1Yz9JUQu311
+YC2jKNM3JD3BF5SyzJ7DnmE4CCZV7hCv1em8V17MeZfvN6SUqIswxsVAe7zGa62
Y533xQ6elDlRBgG6T5zo5I7Zkk8YM/e47wNPQJUR89YDb3dxSD8cukAEMixFNjme
UjK+lHyCCOluT4DErySmqEFcixkFvqZcJZIVlc6eGKJ+mNOy44VzXCJqgtRiGo5f
Hp10tVktZyN+vRTkydxlgopSGbt8sunH0gcyZC5ovN09lQTIrRAk5XbbmPVtr7ur
vHT0CK/UCT2GGzhl94ot9Wk1TJZSpB3uqbvvSsPRiBVdFOyd2DjkiMytxKZuwFK2
+vcPen2H2Vl817duQlSuHQG5ygS4ZOgXkO+k8zWPT9XhQSEYlmJotcpEdiFOSo0R
OGUJK2xHFEbK9nEfYyIyhjl/f+B0zXWBQk6Idgv2VukEkpf1Xz/WaFkBboa9E2O+
zzkftG2OMqgoP+IIIbIdrOPzSHZiyoaQKJZxMwcx7CA38t7rYgYIBXgvR8jNyah5
YSvtwbaH5L4v3TP3Kkpx8wgJzR9MTHCTkvGP0El0DnwaOBj4xyTFKWVj8iPxmvmU
Mh5eFxRpz7KKygeDcs2DBZInPXehR0GO0S4kWsXSmXWHJ5HjGpvynN0pF8KbcnIU
xB8BVWWkEfzccEcaLGt5woAMz+Oemt6bfNYJJSAfnwMhgFXUFrtn9aoVh9gUdOys
ZOD60tLXetiv4jjKSdzr5W7mKNdrhgCdFKw+WH2fUpbNLFJVgvdauFv9YH2t8tPM
rqyg85cfYCXFLsWqPidY+nVt4Aqaq+n5oW3F0FN4jV8Af6RrSzi2QC1vWbDw5KLV
dsArihcQcHbcSVaIQ0SFOXgfxS/cbJ4f52jaeMc9Erdkx1pHMthoOVBmMRjuPmd9
TsguS03YY6TDMKWJsyNse4PJn5GQgPnoKRbY3pbhhjNlgDJ8I93LpbHgDhArR/ZV
QE/maCuEuHPKFtAumVRY8i7YCyLa7NH+F/p6c8hd+AL9Tzuea7XffBIXnt5Q/hXZ
vnjFtIUj/4Fevqi2Jjg/ZdUagzDKaWu30U1OqqO3hRoVsttNbv4L+QvRp+3+SkQ/
VHj0ZvzRKuooUeTB1RHteEF+6HFeQP8jCjw4ELPxaJV0ZJM4KnhAFgwfoGmVFocF
fH2y1+6S8HP0ECC+CoaE85mr3UoYwHEeLYXTQ3GfPoe+0hxllz36Po/RB7eVvnV0
WA3HGxZrJW57zFh1B/MxmO4RAj1W0L1zRc3hmZGkutcad+i4FQExDx/snl5lYqmB
XKH6L171AAfroNrL8YQlUUTHMvR9MLb38CTBa5jCMCuzXZqSxcAZMURfh627jQu7
DuSj4ypEcTVFZa2q3rZ0rDshP5XpUCg9ERzl+Wghxr5dxCU2BCeVlRG7uj/E4akg
TYbBwFLaAMFO1kdN8jBjVB5b8nRMcvhLaxtgMUVP1p43pICFyt+k/Rew0Hw/EU+s
gv9gyUUeoiQy+4rOGUXFcVbvmnkZldvRHNgpVly0700XvbcEcxblGEJq7cpD2nAh
ID0GShkflID9Is3TL/r3t0YPdjdSyOLtCk3bldclS4KyoB0bD670EDktCZCavHUf
E/6Gvo83AuV5boJEcdIUb5QanP2yBiFfIlDc6YwOyGeIlWZ4ncTVd8oSFPP6lYNX
HaLVnkh3MZKZF+rjT9uXYUMco3thWSjHNm7nzRJ/7tuZa43zEYAey43NpFyTm+TL
XEA4FMp0ENxpwuhwFbwHS9n+a6/Y6LUnjlk9EYmYCZfSY7HiHwfJ6ZrT/MKVK1H4
eisqsJ9Yrebp0xh5WvC/JPB7N+wDWSeZBzeQLHvYsGkJwMcSXh3bY0Ahj3hXVOAL
Y7vIg5JmI+t0JUiGRP/k/eYfl2Wv+7UUmIO9Dn2ctmKdnlVH/7Sl717oeMwaS0Vq
ZxopB191u2aAqlaslOslax2I4WtbXdr+cdvFY4a6ouXu7kSGzdNq7Wv1R59yuuGf
9TzyunA3lcLKQhpM77010BFCLoE0YICAOK2deW+7MZ7xDRkaQKFgDJlNOY9eFunU
1zECu6dlO6mThHlxGI0848dg9m6LXjSwtPtYt46/62Hw7aCgvxe5GdxgxXk2ETTS
gr11fqYcczV4ceUWHxRqQGBDN/Ap2F/5xg/GdpMCCEsa02rB0WmLL5Y7pjGk1/Gz
d9Vwk9MC47R3WaGEQg2n6eK6VAT6fGKUlomlkWQHvOByJcst4RflfqjxDAEbvFcG
cZHMln3PMcDv+PhPYZllKFZscDw/06alW09cUZxjQWWoDxJfK2vm6uBESgV/Foh4
RC1YIeHqXtIzfzjeKc39HlO9T+aQcO6yFwj/EX34LaC5l2ZzM/nB9itlJOtKvYcS
l+DD6k75ezn2WcnbSTdK1aesHBaHKF+7hebcqSL2JD89s0tLqFY0wrmLZt2qSOPV
PElflDNMlzkavdpFTcLwN3em4fqxApTq4rxrrXsU7NFCTXX+Cv4+4CqoHhlbhRHb
Pt756fgN3/RG6iLQ57vfmEEFbRS0QQhQLq9MrPOJT2vmmcEFp5hCMm+9byq4LtQz
UTxeCBjgEmDObCAFOZqmpiZWjhxnc8nyO5ryAAlSRxhQTR2ATjBxbMGeXHqK46c+
349bKVqgucjF4/Vqb4xxN+WtjNoSp24+tSVFbb3xOIPxe5kW9kgHMpHMMMujYK0H
zOX0JABejutQhGMLImIgr0hlan7HNSmNobmK/HybCZgjBWDf/96fLrsofMWFWEui
tvMozjY/nAmkUMRWrLZfM3E5FYY8AurUIbbrqoGXYe1Y0pbL+PPp4NhXkShsADw+
8zfs/dWEb3qMo+qHWs/49Tx7YituKyAhznzSfAi3xCg0u8f0FPuLAvuD/BV3tKj4
szkgF6FkX+yV4qd89P6U9Rn0DMwf7rg4SWLcrJTgMOHLG06qAT9gGWZ2PW3Sfn0z
poaN/6XcG6PBpt+5cDq08FU+Agmhbc75OrICtaUkUesOw1sqIRnO517DoNcQ5ECx
vxqk4Dsj0o81IbGfvhzGq6W3timI9sWgWKpxSEya5M1wALxAeaG2b1JvN+jhvN66
irjcoEGPRIrN9K/rcU4Mw8eNmcqLwufYt0/zVXeIch1KGmwjeHNeR3heMp7BL2UA
VdXANJ4FErh1gLcZaRKFezYIPnUHGUobMPby3mvGlxunzWSiRvrsIPQBCd20CdCw
O4NJ47wRxOebZNBNkSluP/NRrgFj9/ehwRtXnSssdvR7vGod8dwIdWzlwSyg5Qe7
kPp4oPnTMt1wcUoTQL/qbNS2cR5p9PDpiG5naTfUP841LaaDntl2G2O2OVsKlmFJ
TL9ydFX59pja3ScDskEPEnWSjaCTh9KL8zHAf7yu3FobbeTC8pr2znin64CTBhSj
xTdvMLWn/6MICm1po3kJbUIyOsAW5XmhivYl+m91AnKYZczWQ2rAHRWU8rzVlYUb
KkZo3zcAghXZlsxbFPFpbytzYu8ZnWnWyZTPY47IX5pXBvC2ej2FA2/zhSw6/6S/
rh1Ma2Mwb1VO/vLWrgOZVsmhOWkbrHxPx2wqGm3Q/ywWZ4FmYfpDvrLuH/wIAfkF
XkJQT/G+a25ehmxWUnMSN19AFq13Kl03yFGL0I0L/wFZbeUmkNWX5nLYy/fc7EuV
WuOpz8tUYYWZELuIVBfWXLh2VXxo0B5nrh85wsFZH4dAfZNtUSrvbWnRlYEsAS0e
5BPOoRxByM22ZzAxwpCigC79kUFaVgb/gar0avQNL7ptw0RV/KobzAkCMaH8Gf+a
fZQ01UuDi/A7L74Sra+rfZu2/DULNDS03k+f3yFIiHy3UIn4z0avHnZpPjLaY/Ei
pKGoo6xUmufrzqEKoqnn1052DJBgNm3Usc7tLZiQ60B07ICHKhctexpGL29RqI3h
3L4kj8zE3mPa4W2DT/gBtREmaSeOCmGb5pnftR1oGVlBdKGtmEE50x/AHQfcTafe
UUAUOKOzVfpYYQjK3pFfiVkZV79GUjw19l9cnNNyIp23jglapa5uEVszfkRjAjVe
+PMUbJZNJKecbhie92IrjEy87wntTUA7DdDHk+BZKYBq8gl9wXx5aeYbB63siQms
rffern34S22UdYoPUO4ECpVubgLEP1ep49FXU2DFgOITxTgw30WajGLuYoLTudtQ
XEffwWy5U3j26ZTAD7F1yVJkPSgKQkRFkKo/leymCJ/YGw9/wpVTN/ue666LPoHd
8xZNmXG82OR+id47dUZySQoyo7jJrzMqOm59sJeNTuDNRN3BcBzb1Eim8ah1Xr3M
A2aqgGh3Ghs8j+4OJLe0bQNlhBIGw/pOPiAELRcVqLi+vPiWpqWMNGfS3cUZjJ6j
IjAjOMOUfXMtvkIwxbmNJu9K3S1WdZvWgB4dhKpYO4zg084AWSaQ0CGtnqHFr+Nb
Nym295XDwpfI/txgHRsk6lZR8nhnNQg7fDrbgJKh5dOK1M25yuwalvhghm1sFIp6
6NbGJchXSoNSdIpBV1F15/2hhJI6p/Gfs8ILjeruX542OxdQpzhJfxSdSqy3RWqk
SOdrWoIWpfTT2OZWxgKkfu3zmxUcS+X14k+bfs47Ks2GxlmkmdmKjywdK53kpaAa
X9BADb007Bu+L0uhDnwmrtEO4g/xRIKiGUVWsEclBCvL2q1kEvApU3/CpjQ8/vSJ
cPWOoRlgI/L0CGeSPN1pOX3G2nzBclnrh+6+RtpIOBdCx0Rm48gmMIpvYBaLLha1
e2Ia9tO1cOIQZLoZ2853pD7py+C5Tqp3YzP6wMWT/hUVOYtD2C3i0pEiqlV0JqjW
8cejfpeVVJrHiXcNeAXNRGrLTxSLA1hkjubLYAXOY4C2e79T25Al9rM3Z1H9CanY
Ukt0iX4a2k6jyju450lgn9KFycf8QPiX90+v9XoJNwr6gKMjK0qY/UN4+nPZ21JB
VwfcAK6tCnHfOwue8ZU4cNd1M+uGM8IpXzWpgaubMk1JQpjRTtWrrgDvPE6YX4v5
rfEq1khwNvF/kGuSJ1yjoAmMwWSA/OH1u1PBxjRhWq+SzDPVMSB6lTGrEw06BlT0
MMaKDOiPobCq1h2JNyg2Cf0EixLkFaZiwpDN++u7eTPiMc+0x3jRTOIAT6SZCdbn
tkejelAnzExLlkR7lsGVPKlFi6r4lAHAeB1IWdqsYFodA4J0soi90k1tZQRWZ06y
4VAEHsCKqXOOGT1yrOE1orO7M9tdxpkxGcsicO+Giiu/+GNucsltxbgyQKMeXVp8
lcNFkxxw9aGhphtGBCgncv8n6jpKzpYa6ETgYjTPAbnZb7NrguGq0qgdMhrPUTiY
qsRQOotbbdOjXB5FPcv88jgiFzRrr57MG5jJ4xNi96+xiUx5B9BQjpB5NwV3Nlwd
ShuQ+DKtXJ/nvCENE+sSSNs1u5ZQ6nnG29EZeAHC5uTfYcmXPpGSYawpYwyHQHZp
FK/MJ6ZzVwrL3LG0/Pxe88maQpTdKMaPDpq3XENWpCFqmlFBVa2hJtw0m6ZMOXu7
wpVBvxpsLw08lRqaWhXw7cRqrI4E03WTFZ5crSBBQrQjOdMoG4u724R/LABk0CCR
ixB7HG+RorlPhcL1eJNqt24VxtylHG/HPU92iRUk32q8LbdXLxUXuHt3ylcwazGa
SHBZIpLCGBvTnChYaiqWKX9y7Og9JsAUzWMaQFqy3UEODTow++FB/nnrPVSkrrFP
UovniAs58besMIyWKlb/ANuokSmb9TFTnXYWVAm0I12yjVakz0hd+zUiTCOc12Pu
UJJe9164xnximQlEF6VUikjD4dj9y6xY23JB7ak9n43XjRKy9NURRE6CRN/MXJU+
dQPEVIUNGDRL0t5yY8gGHX+pmuTv5zT4gLtMl46dypVC0c6waLg1cX87r/J9bQoW
p2jz17TtWTdja0mSMPvJnmN0y6slmy956XgwdjghsWoiftmyKOQxB6zFIZ9OoaNR
QlsoT033TyTdt69sRTy07Ifeh/6k8Loal0HmmFMlJXmXdVEBgD7e7fXHJ0opw+CF
N2mG0WW1jZwY2gUGUp37RARj1gWf4H0/A5MTfzHLL/j0e3XGAcRjQrerccMUQ87L
3V9bto6HJkLzkPnJGCI5Rwk1VCAW9CK3VQcS1zC7ut08fmXzR55JBR1bC4BZzffI
7dXze6hA4KRG7bGF7q9ggkxBomeAyfcds77NoGBuG7hVb287J0hwqgEg7ncvW6XW
b6R76UF/3m/YKUeocz1hs9cHlqLhjUFXDH3b3YpqcBNplqVb6V+MbHHLhjw37eLS
+iXPxtNVsHkoXZbnI8OnuzcYHLAOdEK0vy3EgxM/7WOzUm+jdC2zBr5DEJY6/OYV
+9/nFNDOcfoAx6n5c7Asgw3DXvo/1NJm+8+gIcohWNpD9W10mMybQ7+vcQQuAnX5
yYZUoLgcoi+mRKnzYk3QSS9557kztHN7B8VDeRbiWlW2gLarv4xKvPTCQ5cCIowV
+C2GFWpg32xIJfsN5d5L4+leCTdYWUTTJeXFKuYQspMXhXXcD4CfCFvjCBV22UiB
ydNSdntdRUP4OZ5zWMhZOKfZUO5S9/CCSUpbnZCKXPI1iqLWwtLgMMV09ujwzH4h
QJuI/z6A4U5lrNb/0sFk73WpRs0/GhtcUa/EhYNsZEG8c473UNOqTJltohU5R1dx
RiWbaxZhga9aWBt8TUHJQMPYDFV4bbG6S8FFrgiMHUjzH1xI1Y5EZ9g5+a0htWX6
rbAKM0//vm7TR+QB3GT9sSIL8MaoGnco2AMMcEzDOSJ0mKdHmjA8nv9cOMk4DGAZ
mPaIr0E1CENTLMghU2V4+Htda0equxf7NrbbTxJEC1evG1SKCuarkT3PM6YVI5UY
Ce1FJGbXYU51wafYbSdiSk0jIS4dvMVVY1YT+l0loLWyXzbu4J8cabBh+FG4a8jZ
UaPXlysi26NG7BbwRvTuwbSpimmRM8RuxwjjZ3Pi64950jaWFvcQEsG7Bdz2QRe+
dgTlSJbD3KcF65GryRYKr9uKBA0z+uQHXu0jcDeo2q8Mb6ZQkkdRdHYpG5JP7dmU
Hekn9czAP4qWyQdCLOqYUUrAq/t9pmzTu9K9qSRIRmPPckbYTkf8tTjrLz1L814p
gacWTQQyobYpQL0X4n517BBbsI/p5dn6raExh84Vmgnm02FEfhJ+GzdX2xE8mt84
ZUbozKErHoKbIF6tCu04TOBQMXtCenTulKm61l/sWWMamdeiT5cgzm9IzzgHJuWk
2dvzKrZA6hWeul+L3kC50uC6uFPu+ir1BOyyiULChpk6MiRxnPBoVAdWNwLGMX4K
JQ51LW3cnlPlmfRXW3OSz8mEF+LTWc32PORJFclY88tMb9Nr/tDghECGG107E1lo
Da99MA9Trvt7gUSwaZWoxTajmIF+/B4GR+dHwr1Nk8oIVi7mwVy42KxPV1Hlnhqx
6NZ4ofkpJlw4rLsx3fzRJpNMPyE21ZEru1ZwxWp2zDCKMv+qjXBWemEYb8cmSjC1
XaLyxuT526hmhodrnJ/XX1n2sB1WWv6sNwtx2rFF7s6FMXAa3x2Lk5LdcE483Zxq
fw8G2JPF3Hym4UXDZnsCIBUQR/9lw+M42PbjMnjsb/XFY5DbjS84FC2jfzEg3rHK
MWS93WX3pHmHpTRBUv/8PNJnzl2izAZCod0hXKhmaRZ1DWRqGPKk/Z0CN75go0TD
C/sT+23nZj6peEL5ZrMmHtvmcqVQqI9oNHem96jbsoJ9T6n6+7Yse2M0/j3jAtxo
SS02I+MOcV/9QpbAlKENZ73ms28W0Ym7Ppdw7YEUReLuPitFUxQfDMpNnirnPK52
1IRFp91bHIBYoWdAYUwPHDoiMCEmIXdrChFdiCGCOu2KsSoZwsM/OVWobTOihNmB
aW9I3JcWBE/wDicm/1ioyBQrgmk09x+NCHWQ7iO/zlODvo29q6IA1WonzJW8DI4R
VPTzS8Gb/1SQQHxeXDHdmItQ1Piz47H4aTxXN90N6VJ6hFrEfZqOt5L/XCdLTNtj
mFSe3gKyovybeix1wSPfQ647Y3tOG28Eanqcai+SCdXoo3LmeqNhf9jPhzpJ1TnE
XkEd235KtN5DOKOIsrEj0LIWkIdISuhelK1/r4ksjC7Khk29Q56gxYCRbHyxcA2p
+OH1PcGLPwmzy3pbdSIOHiuKBgSkaIRz01FMT7x6NrlOUmK+Gg3rHMH09J7sw10u
sFrUHDRUpgQXf3pSPcjemdyXsKpZdxolpsOVpzGkj7PrSDFYGE4AxmNEMvmL6kus
nBlGfqTXIdTGSZ+zPy08HgG6AdFx/d/QbjCKBTYoOMcwpIBQ9mDVGYf27vF8gWqy
YiKtsbzqp3pDdjZLM/CxYn80iphuZ5QuThpXudLH/pjHHj2FfImYSa/cppddhV8G
2B2+29HjHxkkE6xjqQahZLwtNT2V5OdMcfqzWjcG1JG9kovoizj3jQg54uXjKFvH
PBzJKiAHmdbvFgh1235eTaGQ4G2DQkMFFPAFgS6QYikGK+JzoCypR/jDBHqVvH3w
KcX+FjFJkPb5DdK1z/MA4sgffzFD72K3vnhUCi6GOz140kT0yMRhrB72bWIEiwJV
n2Wzc4zSSi33VNgujeeZbCtnEtqofvtMRbuC7yG7kBkg3lJGVDNkw+YYAhsfqU8P
3o2yK5fhh1hp3dvsbmo2jVG+aSwZSn+Mv9fsrl8Ua9ZOeDMjTMgkIU6fs+kXW4Jh
3P277Ay7yBnYErCsrm6tlDdJgm3ZkThcc4DDx/AhbCtEkuLqR2F9b6xdoROuDlug
g78v89e3Ldrj4TmSUiGDAkei2yN0iKJ9+d0gSKJzvrQ1bdL86M8G0n7+NMy1oH50
TsxEb1GG7AfiqwWwG9lpRV5Mljpe4QpGOjhs7QJUSm28zEvJWOHJ/PQ/MdZPOFrz
uYvy9lBLzsFF060iEK6xI7nujhbaQHDyY8EkoLUDeZtI1CttegxgVw3I8/59HEDN
Fg1lSwiuC5cufB4SB4t/vxG3Y3o8zsqUKBrLFay8oGIRv8k3UtC46Ik/EDjyvywG
04FjsmMvNn+pJwOzWZhT79iy39QhvzsqB8ZPm8PD2F/MOUEle7offv+6SfgBfNif
z0dpzLsaZIdYE1449JEUKtFXveX9MHaYvawUju7552R57lYBURk2fx2Szk37LhRu
wsiASi019fDYcjeGcl4DK4vu5Za96HFJnPhmVFIF1JzvH9rFS6zZQrSVQTtgviP4
24hR6B0cRSCyDvjCXKQH4g4wu7gVG0ie6K6vxQL6PVLoFLdi87nWK3c4Wi6rcIUT
WXc0PK1vz9sXB9L6+3727lkObnKHs/3oIAl/BE/+AJT34qfc9kvsb1AZYbHyffND
I1I0VZZqZtdilTZ5cLpb1tkYa3B/YYpCIzFDwsPO7M/OXVqaMAZuPS66WKwnJlsr
385PVmghNE3oAKOnQd02TQ+dzmpmr1iUp1gMzOetJXV93vYDnwgRHD7PKtciVFFk
Ngby5CaYFkxMZbzfqtfftNyYCuyR2ZYyfP9/I66UH/Wg1oL8L4B0t4GhZEhPNxcP
raWcdGyj74JhObVA5FtuMEd/eoLQ78jhZX2hp0dHaWKLR8ljS+xtnfbBjKXeyxPv
V8UHzLm0Ba+at/8Mo+uKfGWb9y4zPpgRgMNO/MWNTQQtPpsTbwmSXKqlSkRrFxFp
vsx1WyADVa9VbDukrEOcNj0ey/4sJQ2HxXSzqZTxKuNSojHsHTyYGJpeTytirYti
xBjBYYF8TGW0XMK6+xXeoHnBmlPwuyqLESGU6Lw4hUWQBAGqSpxT4QJ/SX9x7aBG
PqsMJVaCQBfuHhhHU5HqjdLhVuba3jd6+hYj1WyqcU/LBnLVgEAwXKYeKCzGDDuG
/qgByGgVMKvNibdf2gJbo1vtziCA7ywuG8eImcJgFUxldmm3e7se0V8TR0H6gI3T
xFNowoS3Xu6gw3UEbKEDgFaNLXBJTUWU9enW3EdxPqPChBm/CLor+6TQBegtxPpZ
wp6zSj79IVX3hy3osuXuriRa7LJ1/kfMS4KYL3CcfciNbA6yjLK/8AFsJy5UrCEk
gNLVdmsUwWx7g9edTC46j+1gIgecd51hHMyhaXVVxq8DqHS3/OqvXlYtjr10i81W
lW6dF20mRpgkpiA9C3gHiWCam49lQjH1z5E5scWdSXaQRy4ek2j5TiU4rTKbmILY
ITK4dT3rUOUBtbPvkGtKc+G2ff2hxXPOTn/+hZ0WP2KaXU782J2aSfBHDcYgmejF
MgG3JdFebjpuFPuRBPD789M64Lxgvmx3iiz/e7vsK2ZL9priLPRb6g+fezMN8YGG
6m5PGdGe6UISOC7JQXVOopbjMdvs6gKK1/lV0MHfwIwLSnrBtKq8xzndoJmW2l9U
UbbC2pDHsQIUASBKYWi8Ixddi8NDEqwcB9741hj5PXNn2PB4NhORDyn7MiJ9EAL8
ceXPd0QiMeQ3kiavHJjzx3Fx5EmWAR8x3Fo+mI5DZCOQb0eaNpcDGJYat6ErlEUU
DETPoA66uqVxQPmaARxDZ4/uytqOCA56ZxUGmgFBmhGr6i3eGBjdI+TLYeOeBX8h
477BwENf5t0mobMuxsDXsYAFU+ymsvI/maLdJwefJVZOqJSK3sou/5vykWpyARqK
/23NcwqQzpuXTQxoGtlFhc/rZ/J6qk6dMoDm8yy1ynEF1l3A4dcqHtI+y0/rSF+I
DtAEyAOm8o28Vw9o7nfiD4ncOzERBjGW7kwYKqZXNNJ2klhccP6KnIaJvIU8XMCY
ikE0zI/LzxNgJYpCFgf9qjqN19PPljYzL8v7ouQYuqY0j9Q1H627FBPNmVT+aHi+
rEaRGB8qcGej6SRrD9w7EvRVo2WDhf5ysHQZ5XlcCbWhDeR+6DHC9QD/TQobqcZD
/wqTcjaUQbjZ6HhWlx2sDYN+5P6X7RQtUt/i9agKXG8Y4lS3BsSian7YUfQL527q
pv6kYDD6DieGjtsbWumXHNFqeYgDAo0sSk6SY0XJqFHKpkdXJ+QkmmKqUnbPxOZJ
KBz9CJxqYnQLQnupyFnWQ3mKa2cunM8jyw0fNzTTcBmZkoZ8pJXJaE9kQls8aBEf
QoJh0Me/nuQwOnIJANOuk/4QTM28vd51/NIe0A8g8Kv6E0maCa3x7vTAsRrBXUUT
+DQ2QmPbF0Q+B3ZrcveNWo0ebSMh7ro1/zlx0Hu14UI6IfVQghLrwWp2vKoeupZ2
+3p2P8SrFZEzJG372v16Pw75jctgdHQEVVMhhESwX+7D21mlAcVjSlxkboEgPT4r
drw/YRjB7eqmVSysI7dXqHtg1sHo1WQTwSRaeicqxXJ1O0GqaLPMgfyfrY+MAy30
2vEiZ/DMLVdQAKlrv7U6ExEIgMa9hUVYPM7KNIVy+A7lSNp4/u/8HFsH2KxJKaaJ
8kkvXnEhfODx8REie768yoALKt9fdPXHVFV4siKRQbe032mLAot6MFXnUHRfX78n
pi3jhCgkSvvlmd24Qq6Ng0UAm/r89EexPrCBZ9rDc1w1D36bKosSr6wbjzZZVXAs
YxigUF15ltSrzKww0jtswoSx/Gz4JvL3WsBzYlLm5ZYG3b69B/H15zLjkY+vh2iM
2CDOq0EsGXLZHqA2/joTSBj99JPYfo85daktuQfwjJpnpriRcxamaeUs4QMuqpsg
10YltasaXrW0ef4otiaCqdKm3+xDNrJe0JBPD7Xl7/XxfC7ylSnLuHsg/Ydgohyb
fjsxeQcBLBf4+nBI454bbsnRLq6O7HgJ/hOhq2fIHktfOEk6swedWO7CT5syvjeM
iE2TXLwFCnH6bejeO5dlJeDcjP3f7Qhs3ZHRjw1b33bH+v/bakNRaWX89TodEOLc
mWGQUrEWiM0RhU5L8sK9sN47oEGmy8+wUL9OOFeuEVRHTmiv5BRLQ1CZw/rqHQ17
FcAMHVdeUPNUcNHYnEKzhr0maGj7MZ/0MPKE92R2X62AAaHqdEHOv+s85Ch5TLG7
JnJLFAdPtFwvw+XIy3471LOdBuTqSdTtzLRQCJUV5G0jPpphvM+MpgfwSolBbaM4
mkxYj+lwqsRFtp9BXwiGriaKPrOfabOVaiaKqA8VljyPOtw7eDIZ6LLG4XQsd8pb
qSlmoshJrlDDZgPip1359zgMWm31vR8OBsGizMR1z+e6NguaeRM+dDpGGu10KwkT
r8JchyLlhdF2MDh+4yH3l01pIEBZPswi2bm8DVXS5YCAspaFLHTdqypq5ie+B6R3
rV6+IMS2hR79W4vt3z0EQAcgznuXDDt3UYqqu3CqkDYtURnH/XXqhCiDRccZk81u
wSEbsO7WFRxfmv/TI3rSbYS3Th5KHt1NPZ4Y40c5UuZ5EcXcEs70P6HZF1hpRuUm
rnPJ+WaPC0TuY3bM97ZjrMf7cKLqNFTHMZy4aubALqtVsLdVBgiJ1xnogK8r0Kka
T0iQMH4l7VxisH3jrijokZkeIcPPRigqtzaB8kJ3+HkDw8hdd7ZCwAZnOwZX09Vj
y2FONFz0ovxfPkA+upxMJPshrDa2Y6vw7MWexVM3bIveYYfqBrYCgfAxp+BzgbDi
SWXoQZFthnxvv6z1HK2UH22gxIFx4UTYl/8nQTqoI5Mtj1lecwpiZLiq4MkxTDX7
plInCXgwS6JoErVQgedN0LsyB1E1FV5SR7WvWvzZpU71rw0TFA4igcPqkTXuYHGG
z5fgj9Xy/WZbRUnu4O4feVSEIr7ANPqQxapPlN0uRKbZMGY1vk+CtttnbJZnHskT
2ImZ+jXU4UFEHlqtpy2mUNpKFvrKWRU4k1cW+p1Ndg3/yWzwP4CF1qHRcZigv5la
z5GUKAtHLMyJdUxBGFkAgFbB571vpLE1t5zxiVS2qYXwxEoYCSATyrhj8TlLMD8M
sFB16mX8oHpRs0ezZf4r2pz/sLnk6TSoj/a43lC4+XXiv+qjKBUO5nRcTvJ3f8d8
nSf7fJoC3DjJIHWiY/+PKXPWVWdH9ibyxlGLs60cN6uUUl+5Cg835Ytd4WOVL7Yp
l3UWUvGeoBedcYDQk5dfZRyoS441Poj7u/e/LHvmNsa/irAtM20np/bCKILfn6nY
u91uOF3BKihEPxFGUBHLIjf4itRnQKqGBzUBBVMBpSNqFp76RI17BQgFnmIknV47
JFmui7C3Qc48iP88RXzq3lYZPwLNF56A6I8upmh8exc+u1XmS3nVw+vpQAIbSRCh
uFNMkYrvuS5ufw/oh985qoSmxPwqaKPhrZ+CrAptzUrylrgH1f8W+59E1kZozkUw
5cI0bDHWl1+L/pEwJc+FJFx7JGKwD92NT1xymz8wwe+b7P0vFZ7BdxuxlPaJfo9r
iSzkLnFaF22Ni4H89SIPbxnIZ9bUbxa+ZH84qGXT1wYY+BmSEjjmtPWDsWGQAoln
pjInJ078K9Qa0VPfElS4FGmL7NpwIZP2No2FP+xSyQyqz1u1WpNl1yZUZVBVj4J+
b6Z133uCZxOaId5lub3D3t+bc70OvmYeZjN/oPWKgk92et4l30JaZf2PvKPR0uYd
lGT/RHz1FLNJfNxAy49eQE/S2Ty3hSgxLLoPlx5NSTqNwlxsGBHtfHpzJ11bQSab
Y0j9ra9maZiObGAaHpb3yMo2NJPObPKRX2MODHpslFqUTjs1k5eRqlxHB33ZIVNm
TuePmo7Syt3gLFXboO3veYSctnl2ddDckvHyEjOQUKay2rOkgc8Rnh3//k9ZFdLd
1y8RSuFpA3raJIzJG28voRrnit2S+0hJH5alIMbs0DQs/7FBOBfGbU0WmgB1i1CN
DNg35d0WwrP35Sfqbr8dKa41rqhsHtsU+Q9JY9TU7cJ9XpEr42KE/OBtVZm02oyQ
FqqjyO5LUfouG3Y65CJSc+K2UD1WjTs3LGGf1a74LVJCQEtteHdntzFenNozw4+e
S903Lit4xTUAZd7IBWIpGV2TFflF1avhiKNsFxbZlexg0KrfiJaYFb3UuD1vljgZ
ldZQWvPPW8+KryCSC0O8Iwenu5fofeojlXwX1Gbs6NTlDyMS9GgeIQfIKV6sIHTO
KfqNSb9dNHzj3KzDWYcIdOQggncdo36ATfsNWs5E/r17pMcOT9ZvEiBVGurTTYSz
Zm4Xuukbh6nbZxnMUhl00mi/gbAmW7f706yzlwn4LL1PbmObRfG9GFs4ZnVjAG5q
qPFxk++iijVxtisQokviJ5KAqSbQEcIpGGUbsCoLYgmJu0Zzw+ejxyo8TLGLqN6Z
I6AHcStfWmNc6I5brB+iK4ll5IIu1mvIP021WVjQ8Jl73XF76E2o5vIVpkP28FOv
3xkW6y3T4XytbgHTgD62DqPvnK81PxJfFd/9wz3icLjnkXyLD1nMoTFFOlU9RSn2
ZiNTKwLCZXjwzCQdHkM7lxN+xpEdqMpHkyhM5eIFtNpex5qdNftNMfk7mVQxkG/1
k8b1QLvcBL7Evr3aE2CIXe9m/NuvLwZI+ZD/dw9SdBa2Xj2BV5EdsAnI30AAzZ7t
odulVapxdtF60sw0WsXrCwbscat7wKw7dUBDkJvOVrZcqWxeeP2vUjE66FSyZtcf
VVGWAqsuBwbmN6x4Pd++WAPJqBnu9HPhd0QQSIybKrvwQH2+jpk7S+Yw+VcrTsaT
qzOFm8yZ4cY6tIS34rE881I5Qacz8f+8ZyC+SiBDe89QJCEkijahKaQP1UXVzYDL
gnXSpmrEM/F3odk+SwJSWceaNLfjwZX2eLmtnicabrUb8k7ZhM2VxIuVZVZJIMUh
7CZeZj+Up7woDk5zk2tiUnBM41SidgkcZg5bfp2TDSo3Dt/4CWRCE0EAar1ymoIt
X+86slefYVd1ZNeBRDBbJ/+24vRPrdg0W+nmVVCoHLHTSDfxNhUG72VFPiWy1LHV
CrML3u0crYblH506D/AW2nFruBWxJMn+pIOWJEmBETmMFmFyOjY+dSLkBgrdiJiH
/cPg2bm3eaq6Jk/kOXtb69rLTNohVGSy9U4LoBBoNiRxYNMtQjbyz5YVnCHcIO1z
4t7pLkX6kuZykuklc68Gwy6QoshbVQ5J/4ERnssV34I6y9kbHtqbEQ/JOH1/Top0
fU1h9lkFqMix5XNLtJw3kFbnT2Q9b0c5qUigFZs7ZN3qGY10PI6PhwdUrv7whMYS
6NkPF4+HxRsA42RgU83/fai/xdZu/M5aII03aChBqK/5aQcG6h+W06O/VGiysM4h
bs5DGcaNkgEV0x0AD1Zu/h9N/TEKX0yJaXNX4SCltQuhu/p8WfBbJ/0utnCjEumu
S4M3oZiBhjrzl8hrFTB8E7+loqPJJYXp3YdTP9x7Aa0nxWTg8RDG1OR1iU0/h2Ce
PBNnDEFUKRnPWMhm+iWsGUT/y76oDpTezsMF/ZyzQ9EmbBJ7nF4QhEn5FZkefUzt
jpaqXfLvvMz5D5qqB6ZWaUR+mLFg9E88Y/CKuggq0Q/k7LsaVW1FZdZBcCPISSyH
B0oKHH+lkHxKE2ll6ljRyq7z5pbK5V499ysaGCAdV6V6VHdWaH0OD6cBN1DQHqOH
+CqLKCEmirB8kERlD8jv76lbieIyEr47U+pmwgUUrU/rHUj99IemrIjOE34Mz3G7
lO9Tma9UA0wINzlxj6sNUQeLEI4gkSjAkyQlALhcmVuE2Vf0M1E5rHc39dcbEVmV
nSACaQPn7d434pxRWdo5FE0xQ74BBHeAK6mCEosl+ceE5z/FKwI1wl0pDbfntqw+
sJcVTv/4urAg3d7zov/K9yaE2pETahWqbevGQ1DXfNnQU6PIAkNdwNvRxfDng96t
BIGMnWbzyDmQ8ZphVv6MegyyesbafqvaigLDFxecSZ6NTeRQoJRVUS81clKYRKo4
fSglSkB9TeJZbBdDEgyuAYh8JUACkz3WBSoNNTNaGM2hhhljg+7z3BWpAnR67H4F
cyxOLQICbwbDiejYf40XGAZIYmHU6jFTJ5plEZkr25xeBfhMrqG+s8g5NofEoJcI
Dta3FncCmPvj/D4nyNSu7DMWUEFNBByHbAgfd3blQD0Ef273LVXeQ4xE9jN6JFPo
xTSL8pg05sagwihh7P/F07Hg5OKK3LettG+XghLjK6fZQbx2a1VaDsPo6VacG/8i
lcxVroaMIcMJqC1j3wKdWqlfqXn+uo+qxzTk8osgBoB1s366SI+llqd0CapZytsY
rpEyA0iFEptuc2aoqRrIk6luy7EyRxyZxoxwBVb41kZpalMyLGBov19WqYQZ4cqB
ayH3lJ3lR8A/L0fohv2zMtNcv45voHStuWf79SdOjLKtmb3/vBeEJKyObsZCZnKK
CGqD5eduI9JYgehevO+Yaf5GpeefMDmOnlEQuNBVpTL/mWh3GBafM8qv7pI9IsRE
dinut5eYuep2aegGwPk9KgmDbkNHdZNyeYi9I0V8R9bFwyRD3yR/0oyS3S+Gn05t
dNhfjKNqN8tlFVikTq66NEmLLy4CJIY4D1kFCxjjrrHGDlTuG+eTY17wIUCx53e3
8O0KHzURHD1S/HA9ugALACPQKOJMT+ZNz8i7zNlViXn9qCEOIxp1k9CFMigVRuv6
9Qw2q9UTx+vnC962sVWBu3jNdBXzhmqgLit6J85WvXBwcipmNgPf/QG81qmih5kt
Zk9NDheFEALN4hKDDZ6tVdo8spi+FZqIQ/547y/aeyN33KfZgR6j0c5UFcFTUXp8
0wOTbfI9Lb4fuEzFYEIOCij/2YfmD7yfxovjnmi1EOmwL6bk34XpSeJDwf+HuYH+
561gVX7qboLXkUlj99saJcg0irHZP214DwcKviXvvFcv1d5Vs6Mrne0NKCQj39sg
9AbLno4mqVRRTXGBKMcVC8pdCtiRgLTW29TwT9CxfU5eCo4lgnWtOEkE2ykYigzB
pGJJgSWFWf+hemUyKAk9ZQVbjlnoumayM3LgXx1ilRDUbD5Ma/m8+QAI9LkrQoxa
qyizLy1j0KINLQTmv2BsOZNeANFphjiSMPyvy57Pe9moEZbrCnCacl7sHsvhtwIa
z45CUWBvOL+M/uLLY/eqTRdSA2n+lTv/9lLdDQoErb0g7f3jXY/ENQelw8Gv8Eyb
BFLjdIlzkDvjwE3Nr3av9B0oFpZB4jpwHw1aL3y8I2+DNJjDEllGN5kvVfxRZZAv
ZEuga/uQ8CwIUFjGofV6jj0xC91Yg90X87sYuMSmZ7H/NQdJ6y6RtBcw5zR05X9e
Pi7gp8X5Lhrsf07/CGdn9syrt9LYwxbijs6OvLg22IcxnwbN+G+7AxUDUFJzzdzW
d95Re7oz4kYMdLONi+GS4rX2I8cLMBss0p3FRX2Vas+iSO4iTygqWAqVJdckpRV3
fAvb2A0+SkXOE68D99AT2HnRCF2v3yz3KglKVbTAxOm6JpVO5GK0tgRlFTNy0KAA
bGAh6A/+IkJW0vvwAlUtSzE9kDXdetuaBNMKtJlTwygj9KBLHaXQ8Rzs+f2JrRee
s+aqgJUBAexNZVkV+u71Gq9bVmhAyhu1Gz1L5jeh5I9Glks2lTzIJOnhNg+KYl6h
AnaYRaJUJRiUUNLYXOnDaIFCSdU/JBVkIfnXV6W3Z0x4SdqJ1jmXMilwQORgVqZg
xKBTF3wRTPaMqQ30bNNAb+Lg/8Iq1MyGAWbZUL5aJjD9jUQPc93hjdzFEJAej7bj
RbfpV7Da4b9uMOvpy1AMgBzcjLK29OclZYG+ODOpGIgTdnJNm//EtHksRXZe2Mfu
Lrmt0OdwpoiM0TnwhWK/qhEGb6PPC80aSSm5ILHIrYMmRAknYgClCJ0LbtqoVfju
LdJCgJWGxAawNsMSS1MATiMV21ETcjIjCZwLu71Rx+/mzG+pn7svg8xJwXwMGjTx
UsygE1hkeZ8vdgioaqxvsIys6EnopGbpsuXHAvoJCsDTOKhK7nP7HiFBZOTE33cG
8gqx8nBsN6cZGUT7BZARjTNy9wxjwZGOykA1LOMdRvW1cMxkbIHpfdXGRHhJIXqV
X7wcPkZd4ZwYvqzbelLL8oXJ9iHQzcmD2YLH9DVsTwJ3KxYMRnD06XYIoH+H6R9d
2fh1m9jEKP2ddHDZMmERt9lI4mQ2nSLikYeXwKbCj46quO8MU8YvGG99WMu/T+l4
3QH2rnxvmJdrxrdcfWgkCtoBDMwDSNxqGdOAqH69v6SFN5h4nkis+NdjSiZye1eO
y5rwYhHmWcdX4TTN+xQqgNmIb3OeTutXQ9AsYbX4LTnrTl4HhCmAsDxjwERxX6NY
SbX9Z52GJVvHR5GIqFDApKLwGg0T3yhjY3VnDYZ1DDa5Yy4zcl1PXuLydnGShuDW
8BZUsFTXd96/q8M05TrE+RK6bh1nB6Guz81jcGyyQTKFvHZK/gYyPnksLE/TOslF
326acPMUeFhOOnnJN42c95LP/F+T3IpLi3tiF2IZWPE9jJdILTNYhMZUoex3RjGb
2MAzSfAKHz+MZ/9JThc9X6YBQtJKqdDvQGyCzxPnU+ea5eeuhbcfsLvHCUIDXLbT
ajY9Yg/m5fKhz+RSWpdCoXDD2v8MdD0O4+QX3eR/IM5N4h6XmaDX2aKNeNSBNtso
ZJsgwtCZ0Tw1J29ujtkZOx/8DeVPgtRLU+rV+KMUDT+hm/MyhpsFTRiVQVZkFAou
RGZrG37h3syFkTkL44uzl9WP6yclof1VBJIQ/88wz4mtk2RFsKjtqEkOlb7VIRFj
KZx2/3E9h1ldRcUnEMqm/HH8QDcfAELaYU/HQgV/zAeh4jjTdzAMAOM5Cy792PfG
yLvpadjGLRuO07lV6ps8PEIvvUAkOwgt0msyMRUmvaFLIQyjtABw/izmKYos0pnW
XPuj7q90ncRNx0CSPmDxOvny+rWlUjbSu5SIB1p57enVdIfUPIcnsyTB4byfeTr3
kCJprInSxAu9PiMU3h0+d9wyyz2WwDqhwYg9F6L2QNn3KnQYscFLISLs9boO7cUb
RY95pB7BIqGZQGp3y8ELyMrQmoyLXNlaaqV2HouzxvUfhRV+Q/vDSG/vvS3ysQjX
Wz1S2zZ7/hdwvQzroVKRIRssb/hbFGRDf2uDFkujAY447agJns5A9QD0ApL0SUQ8
Oe/4skD9wN5ImKG/nYnj3hWIKe5OYUooYdpZ98QvTaHO/wZRqCtLi8YYGitTGn5Q
QafIxEcI2r150h6EEtnUPrxW/1kMUH83cTBAjnrNYUHNTbChPRcT6XKXRGialhcV
Uq0aK3BPst5Za2GOlDn0YE8j4UfLZ9u3BU59WuuEgs7KDHOktsoF/RaDr8eYCD0F
B3mIAw6amLoGv0Fa/bGpT0MZKGJV+F6zFbXBi/ZzDkmPFHiuBWOcm74IWiV9Ju6m
aB1q3qbbSXyW7cJr2ckAIXSFzq36X1RLoSZzJDzYJMkbW5cNrS8EA4iGPpB4VdsX
Z3g7gwRZHPJISTbOl57MiVFLIqibJGI7/74bnvRJzhEDdP1om1tEWM5owRv1YXPe
c5LBMwMhJ0DfN5dbXtchJB0YAuT4ki+7oK5i1K2MR1+EQFJhhsCwnz29vhvbl0jr
/rugJUEDtyYeO6Y0Rr0w6Hil/bi25GJtJeL0F0tLh9j7AvGEE2Bfd5FtHtuPd5GX
ypqFgRAizDsA2QuqGg8Yvwf9S8XbI8Whw55P34LPUwY7QF753Q3d7dDPyAHHFocS
qcyQHL5/lck3qTowEm5o1nAoMyjEHG/WCY2XS6+H7iC5BCvJZEKDhPNluccyvqeu
AxOqySyQA3sm+Rj3nhkfbW8ldRk0T1L1tgWE4FNWcx82wFB1QUHsrOMPotfHkv1c
qQR2JdKFZlwHskXl34EzV4C5uXM/HkOdsXJgJpLbmhg+VzRkkYi2z0kJpW4Un9EV
2ghycIggMV48PdgESsOSF3lGRznj6Pz67USD0EG4jprQkuoa/L6pIBJc2CRNYYEQ
jgzUVdhKRyxUxfhzeep8Mx86ivfNh5RR3M327gO2n06EQp0jNg/DgQSMPmMLgG+B
+XGLVGNJ9dNupkqofpSvpz0u8EhvuEswnVtPa6xpi06BeKN7VTnN2vbF9q2cv6LU
0wKefHfeIVM6Sw7rMKOOzPBM9yQwJCMFOPWeuTvadbrhfu3fxgZRjcQzc+P+UsWm
WD9oj17nubhXcePz7ChGddY4+67EBE/h/OgDFcEASNEQz/3YSBXsroEgvE6bel2g
v+GhE3JPs1z/OfjpdXytQOHQjteuEJfWjFVo+p0Vw//9/ltpVBP8YC5/H/eaW96k
01uuIP9uuQHgwLswTSpMwRJ/sM9o4uPnCpFPiAcgNVM9hY3SV86gvWtCKFlnPIfU
U0+qPweMo+PDlHwV1NBul8E6Z6/136u/2pNJAylPsFqhfUP3+9h7L9J/ORC/nrKy
AFDH7brepQxGqDF7VirrrN6X6gGn1YJHYbkb2mRXuunZgw/6AWOhMr/mnX8HlXMC
Hqq56P2SuUv8jJFDteaW5mTgAyGy6rRshu5NT0dDgqT/Lw0AOqGK4AYhTRMXHB+C
NaoAEXMavpHiQ56MhQ5FP6e53xKmw/ZMbfBl1lppK7yFQFN4njr7TUfKSdPF1xuR
OSHcp0wfISk+zqOZp6/oznJLJbh6ONrmEwa/XLS/DSy8iWmN2Jao7rpruCHXkS0P
+72dk2cmpRsYG4g3DDzDTkzFbLtctolJrLi6azuVUugINYKi0CcLSS0C2CMrcE/k
gWhkfWmEVx/qgeSx+21s/HRxPYtY9IjQRBtGP6LZk2ygHaKT5ypsY0iOVi/9eYSI
nsqE3kswK4nARN6EW4Gk7GtAoMATlrKurRkLPCz9J++MDVrLVfMvK4ndve9wpOuY
dnUysX4pBMHNnzaWN5jarupYLAGgZw05rPh7C44kSTmDIV35t6hQKwy3E7Xg7Car
Hqv/j5UF3ZqKg+P5fu1zd+Y4+9VIhF4lc99+fAKQIZhQ+bZU/jEz13qvCKWzWTgs
wDM1hgIRXU5LxzZSv5OkLstYU/huyAYWwXLQYb7vDp0kVl1r6NzHeJmaxv9LEidn
OGNMFOeNfiHTT/2cRfDYhsuzLpJii93nlIRJY4rsi09HMfkTue+ShFkXoPkhawGe
Aey0u16jdxLwafG1cYC0tnObA8YQ4JYg4x1uQ7rrTiB6b3PL8IwQP8VXjkXK7myX
57zPkrokAX3Kb6XON7Q0gNzMNH4joVyQ5qlbGRFRRTMmG8O0Ugtd4KapcCBzBsxB
pxISj6QBwFusz4qkm7GUHaASGHYa7vF50mSd6U0KpeoJyZcHv7CZaFhtCR+dlrol
kKn9rtHmFSCpO1Y5Axmv+dH9RW340BeQjEF6hsIL9Yv0aZiu+aGL0PMEWH1Uu8GM
LWEdt7mU6C7vh/qL7jStyHzbx4JGmxoLEZZX8Q/XNxwE/LooGRfOXQ9i0K+umrei
5M9pD6Gjgf+Qi63HUIaofosJFu1EwinK2cggDDbxf+O7ogHO+jJBBcZWGadDU89+
+LEL5eCX4qWxGOy2tjlGi9lL1qffwJXn/XSUDB3GoNK12H2IL7t9JIKHaTR1T2aW
qwDGtk/LYMe7DU6Y71kYNI3dvAVbB7B1J8LyPbJJbO2VKU+JZ6Qnb9HlBBJQUZQt
a4rxqH6PBZNjgHsLtd3+adSDu9CQQHjruBiVVRhNNwJ5P30I1juPJ1tRGMzL2FQt
gBepRKewaXqtGX4kG3aGaj9NyhtjD/jnOmAlbxo37ZTG6hn9MAB0/Xmi4ezKa4xg
3rpOEmCHLE2UBiczxKOb7qCku5DGBNcmtS+IoWe7L0E/L/wtx/JdJSEi5WjtulIc
XvMmMoCfsHBzQC+Hc8MQKbv5Oue7JhJK5OKT1BZ/o48ASovDVrsgaEvGI7TRrW6k
t3Pgq1B0iQFPPBD2uMOtv3JuVyodK9qqPTLl3ZrWvipCXASoPub+G8ydFdeYUpo9
g9W0U6zVO+jZpVojazGps7quq6Jpdk7HzyJqpGRbDjk3S3NCZF8Znt5EBNuuI5Gf
E0IUYeD13cGglTjeIoizDmjtjwfDCm1+kMzLxbh9m/byJl0LKrNwQeQUZU/RJLpK
i6Yn06ufOD7jdvV3xHoofL7EooTiW+xew/IpaJBwsF04OCWDJDmJwqPvtVompDsx
43aGVzEH5ZmyEuMtIDZlAQrbaVbXGc/pFTLwfcxnDSYDXAVja1J339WBsd37c5vV
Ym0eyuAcXa18xDT85CRznDAz0AAcCT/hzzeMo+TPsPbqPxPHRPnlF0F7KHC7njyT
hRbwrYue5ZII4wbtRXcPrgQWwWgg80zexlPFv2LZ8IaGQnQQZS4PBAf6KICrEF4t
AX4BU9PnRkydG3AXJZPPp17lteEjBhTqoi8VCzBMGKfWgOf6GpnYSkqPDHzlOe7E
TeoqA7a4FEmB7J1tzwLlYcT3ySek3A7Ct4fO5g4+OJvlM1kQNgwwBAYnZLRw9feh
L2oeLr0AM+KrR2Pu4kpSiHea5mfKl7AD2SJkLt7v2J9+EnBg7Ka9GQU/+klkJK2D
qWAecimpwo6fqxjF0jGDzoJuAXUojMK/kAPPysMB3lZwV/j8UhsqEXGuJy54Evgu
rF9eDW8D4iGajhuUireTJbWKHhwqKQD8MseijIngkxys0rd2LPkg6A4sHD2bzYaU
/VZzFRzUXVUZouGLC8hCXI+TVkHP4XR37AOUdBoZPH1AHu8evjScBLqI434MGuIR
SJPl5QmelN4Bkp8Xy0UoRX4bkbB/TqdEjb4jQnzbjlplKAb4sp9Oku/ZRtaJSGI/
IRHiVwcnAG+T8yEr8FDnx/x9SlbQ0SYbBipzDVFaQW+CRmaMz9TcY5nISQpkLOqO
JoaR8SyZ960xTwdJmRSfQpJgmyrubn8jnfLvQHt4vv8ba7rx/ER9E8DYSp08hBK6
a3C2mxo3ezGNlHBkTMo9AmRjJblseOhH68JGjz1nYrjcA4PFZRjC3DtAAt7elYdh
X6OH5itdXzjijG/o5ulmdEuRurkQCT50TArbMhzjcFOAE4fQKTQpxOxPYWAqc1xi
9RV8BU0DwHBxB7yWVtz4CKymwfD/R5RBkKD29AX0QIUk/+I6t4gS/r3UzaLXgjLm
lcnrGjeOLcaM9GjrbVc6usbQSCRVOmh7zQXKE8HHbwMknZARF31I16z2poTrLPXD
mg7H/0fHgWTgr6JmxIfbp5Z2K1p5fY/CtT0WiwGJY2qSh2bYpi5rEDleJCUd+oUT
6obZV97/tofAaIcvRDI8/8oh/4K9W7AtXktl5AVmZVEs+tLeuXMR3VZl5do3pktK
ObnDOBdw3dMaMLHJdKzKKsxWeVGJ93mP+tVeXaa7wOtU0ZbvQOgQt6MFOo5Z3Tne
B5fG5WjBS2QT4jAeieUBdsGwfpH1Dd0EOhbVsjE8N3hsnzW4NoRLHQkAs+OLar85
MA8Ehifudjz5Y6eearnoEHwGxtkGRKVjNDZKdjK5bYwi1DrhAMW1QxUuhl5SlWLd
5gpaS/VBpWPdC0M3ZvLumC3zX2wLKIs4yY0T366wPoZF3UfvRT2Hg3UHcPhsAUyk
yeVjwoq+GdFzZFetPtkGTNDb7CrJU2AovvVzMqozCxdIJ0hHeAJZqhTkSqxnxK+y
0sG+Ce6lzUwjCaYJakKKmjTrCn1VjHUun7gberksZsjoAY+Nox18onl3o8IV2ptK
5+ss8loh0qPg1ROEF1Ern4ge52VuxOhvUR/2jvP01GSrjAWEmbCA6rUZ4PZxp5Z9
ucbZtjH8t9gMjZxy5mVlo6xHqH7NggySxLFgcaq5nPvrIUvEd07mrOkDqZAkY8EH
vdnBkzriLlgpQYONgcYftcjyuHQhS2N4nB5h9UW6nC3LJHTQ8soq8F2cB2EEfHjO
1UJHN6AeUplSWnlTS1v/k9fWnXzXibKVgRlZ34Ol6IxGCpTlP34eip+VZPoUKc30
EL6sS/ohujX8GQheUZbbBMZV2bC45E4Mw+Y/fEFxLgZhzYIHrLswwKBpOMDHtajV
5WZSCppgksYfJsOJRLk7XlIQUUJhDPVEUPlmMrw8HebMge99pAMDjOoeRPLLpG8y
FlkFMbgL4SBZs+IzBlCk29QJai/0xPI6lFCEvMgiWprHqiAj9Ctfa6EdBOL/Ppi1
H5hTOapeLevXx89AO/AzQH/pOaQaYNqvZePeih+vmMYCA60RQEBCHz9oHADiODWA
kFwoenZxGuPF67uCApwAmW2bUqrmu/ZkguqBcKnk6ClTQhN5vxCHpbHRYtAPfCgX
hN8IV3RXZJGT4eL/TdFqS0zkgbBEaRkY7S13O4EFs/+BnDANT4ks4X9+CJ3eMZ5g
DdKjFlmgbDRI3aZAbJ43SRl1ia0ouXVzSUEosIXDni1Pq1UJc9eKmuXVRw3msFq2
9OgBlXrWl79mzxs77fF9o+ZVF+AICcfVvQYpX0vmz2qCCUujIyXCwZyxVFXDR0KI
3i2edKprpFH+G3EKSrg08GeK71LlpHy1Rs+E4J5N84gFLCQwVw3MTqbobhqOH6Uv
n7mItB/YpxM5le/wekock1CzQ281i3xgkfDhERQ8+LYEV5jpBcPFvPDRrs+pI56Y
o6WkKp0Dg37l+oU1WnCgB/49d4tpK9KDxZbTwQsqVwEki1VZjYnJQYD3cFvfjm85
Lt/us4UztEpmI5gHmxoKsxzGz4FayrVZ9B2gesEfaSIUCc0m3rMgu3R8IYb2AQlI
Ax5kbycOPitZ/9AL56EAPO0sUOfRAuodA2H2F/H/4UcDkg+tQ0Z+F3Eu8D/wSQEj
mXvmgMGzSGjAuG1l/MeSNk8br8BfHoP0vF2poP3tGhBOIo71x2xPV+wV63AUzT+T
dGUWmCW3tS6YGeqWNhg+9CBqPqP+VgBVLIgImNvSqPGuybMgXYBOzWVc5jxvqIpv
2bjk5jBPjt46dQosM5zK0CeYMzpb0SG05x0sAJuOAjDGY41Mi+JwIyVuS8BYT/Ul
1TJQEtaqedv+v+7NY6rSLRyh8xcuaMzatr7yJLiyEGMcOhoiJ7y/BhwmtbLeEfZ6
FAky/WnsjZg+/PIDQq7LLAd9Y9H8IcueiFK66hOcd9R9bKi3UM1UlcS7ioxvFEbj
p+X4d4psfWhjg4bYRAFTOxpgRuIYBjv1+R0YaXv436U6Y8XjLlADgjOqEn0IDUzz
mH1lCQPcLEp9pxmVI1clAdhObTWgN0a61RSPuj0sg9g0MS35TvNy3+p4E7StreRL
2CSozL/J/Ml0AO3pbSM5flEVyqtW10Q+J8sYvJRiMmVMZSBkRQh97yI8D6M29YML
Y+h1nKh+uIY0zFo5/yk5VlpwzroxYijkTf+h5KQxLw8BumxJ/vDRtBe2NiXqtd0f
pjXrtjYaMRuh90hKKGty8E43sVGwKO73lnFFweWgvhIFffvl/5s7GFADa+0loxuu
rA3XhN17Jihn9fZx7PT3OjqShFobiS3fSqmOscSInAjBSnnMA4VTeRVCwmRBOOx+
RxEZWjInTpdQoVNM7PoBl5ksCWea1ckBKT0BhjIcMVxlxGYk0JvWrnKhFjzgFaIJ
L5vFvOq4jLaab/3GZUw2zWlgAl2JKzax2WOOf53xrDSkNd6TKOkIma+JEwRMEzWD
I8ers8wFJP3+AxApRQ+Y8MD6FafCGPnvjb/6gIbFyxjtAmoFVsBzEUBlK/nBF/Jl
K3p2KxwOsuZMmrHZ7C8eFPn2BfoiH+xrTn+OaeDZiabpzWKMJlg4c8Dchs+yfvyl
U+WOnzmouzA+OVnDZleShgITE4SS57g8ZswWQwxfz59zsIqGLkkhRfywy2T8fEML
2WRlr8jTWN8s8e/ePdIwos0panWTN+zuF0edGws78gax6zmgc6cgJMM4Y+Xx1VOq
AkmrKXZNGjJ8iK9t6UMmCdTJ4rPDKmcA0D+gWv7T6t2e94ulKLUekHLdZDSnGPYI
ekiASfpG5+tAUSILjpUZbsVSzBONyRezLYjwCSbjE3MdoTCeyk/nC2l37358UU1c
FJ/0ufjKNzh+A9wYqxbAzsTuNgu40w9AlSTxrIiLeBLuNgN4npmckeGrpyP4Zu2P
lBcX5ZqLLAl5S1alpsIkfH/gJlVXrGBKtlGVVln5Qkicr/zSN9Ch8llEt4HSi7DW
JZCJil7bp93UcoAl+NvSVO5QLapXmqJUHLRMHJuy36UyRbrXe1cgMNfP+Xpfp32y
eETTbvx9h1E82ZfpzIRgC9qV84aG/x3utMzxAa/2KC++sY8vwaD/UiqqbuyW4kHD
im4Xn2ybsfvwAl+ryC3lr7OfhJOfzstTPT0QjAjFjnOqj5YJsevur7xehy7S4YV5
+Sip3Md4BJr3xJbzjue7FuPCtEclpL+UKV6V9s2Qa1u4YtJV1iGltbBUIpaWWyUT
dea+AzXFDHfcDuWo+Cses/fYMKuV0X4ATdWwfOF/GhPuLBVkp1lFejWX9zEmh7vN
Jbxg4kfgZo0aEknR5qsxfVC1XHsN7C5KRg9zdvHLuNmnn0gyHBbAlgRJ65Oy+kWV
zow2viZtot26XQDBJQGlElEBsdx4/24sx5aZKMVsBFoPphS4r8U6T0uYUAd8sxXp
OAxV4dN2baIkEIZBNI0apmtShi6n2th/0dyyBu83wKIYhX1IyWxu/vJW2qUv1wF3
hkJKfoQkd/cicR7UEDteWuZfLIxD5wfEg9p2R2OMMQTl4aSsG9FmetshcN6HtCX/
PWbj8y3ZamEn2L4g8hjYlRK7YQN/y9+Xvfb9zwr4HmKWXPcScf3FQ4TKdAN1XsEx
yDwbOnFGYkjte14sIDW+gmgXYJYNhb92lt6BmikExS32eqJC4oW0jAqz+56BlISN
O863V8mXwmc8rzfmVKpLWNJGcq7b0eVQcFmQjrG8nMOdwd+BTpdJibYXUNoah0TE
VMKkdEA15WnV0LFJYvUx4zt7oG6OVtmBDiO0xFujxNFF+lXpijwwYZByy6QIZZYf
Bwx3N97NHama1tpKrDyXEv8YEtC80ihYhUmj5USiIcvRozObfei+SuT9x8ljoOcD
3jbZlkQDrZbEySvLWmJvpM2zxrs1+CTd+zRCMZqtAF1bJFFju+EvlPhuZlrUXmQe
lf2Xo3Uv3yK9qTK/76/ImyW1H/CWBwXdTI7bWQjYUo+tPrX61n/YxZovZAqjADK3
egST7q9fimts9GV0VBD3PjQICnrdSQ0uQvboCdHmGI3wpnWTfeZNu3k1g3JHwJtu
v/sdcP+OppXJNG7bgfeAwgFuh/nXzOBO7KJfT9klle7OfvwLyIQv/AOxNfHR+p22
TonRKz6v+ApgY/G+eua3GLuInJQ+X8NPe/T5yoIy8rjGpBN+V8BxzIlwX9yv/QOv
uXlx5wyUrBjT2AfKb8i4ApW5R2Vj22Di1Q5FLtZnU4ajg+PJG2ZHbQUSl634TM3F
U9GLU3521dGRTK/NFUX36h+eYJMA97WG2aOY4i718FCwgLhoS7sRekZIkj4x5tir
FLGyOTmXT/iSgNdxKATamRjRR/7d2EcZK1Fmn4J49qyOt3nrTquv1+mNl1AU8UJS
WN+6ig83pOZlKi6jnQKxIHeK8pn2AYnH5YvlXjPILNnYV2QgsVgmEof1Zuhwf3/x
9VBmLrIEOg7g0/qDIV/rI77Sud8Sk6turWBs78SiQnhCkwPUaTjs4nejP9ISZxSV
RdDL5CP8jYVM2B8k3WYrP3Prwc0KvD3P568ewlWMQ0YJN0DvmbXqs8doNjKNVIr1
WWSA+qSVSwgp8GWUPTJpq2UG4B/zQBw0WXWxc83vgSZFip8J4y2lAK1X6Gkc3/8c
4pGuo48l8n+2p1ZOndartcFkriQhaGOPdvCWLI6M1CUlP52PAenHPTK9JuS5/DV1
9hJfVo/UzEwB2VCxJDus8wCoNqfxEb9aOFkM5vV52jU60yyHzay6JCxtdlnGM5C2
JFQG2qHbcPJKmoY4luYe4nAYdlO3n3gGIzaTWzghHvNLNDXq31BTTbW4yTFIwIcI
dmgvSOIGbkWJzBsP3uTHWvhOgwKZ7tII6tThzp8PlQoxxVZhuWMCiHsdvpOz2HXI
Bf8sx/suo43CR2d67slwevXCmEcFLrCwFDB4zxDoyqboeB7HBDVLw7t2C7SIvvM/
b3GN+Z218s+d12yqS7Cjy0OKkIy8rDP4+UF7o5caRt0N9VYNyhEl4IFjBqlacJDN
1OkaBopxJ+pL2QZKdv15vDvyHR0jhMhx9JEcClWwjItHxSWgVSvRni+kRz5agMTN
ezTTA+h4Sm59f3qAjkKd+m2JarKk0DTgu/kESjhkRZwE/AYa4stFD5MG4ROd7/41
rOBwKSZdGtnuRL5dVZkM2yX9qqRFp2uxXxUKd6UPwylxEGEvfCEuTlQzuq6U4k29
O0zgE+I3Jjh42+L/2HB+hiRiILCvWL2NdBYquGgVATo1uOT/LHgmhNzxf9k/lGiq
D6Ndoo2Md0g0aVYTAe1/CDvGLTDyS6H/ZaNYYQ5uijGi0FbkiRPWsn+o9YXS4dHe
LgQkxwCst5m3tIdoogOXuqdTS8nWOEAd42nNGq8b/0foSxEuJLGKa+YuIJPkF+lR
F74vshSmAAbbQiQxpxDLpsK43gYuByHHhWpXLqCJKujkjfV6AIRfM0ugJwSZbITU
Dk2vCgmwscASmGE/mGqmt0bLYUbXS+uYsq8byOZFUd94nQmqKLw7VzG5wwrmm46f
Xjk60A/RiVuCjPnWgkrQnQFT4rseQe9lh9HV210ApuuVHxK70lIilSeKh/RyoigC
veFCfr5XDmWdnQPEAh4SVoA5148q08HqFxzl692w9JbgNKSrlq6eJ9Zz5k394fRP
JOA9uoFWhqDc60qEEV90x5D8pjCNM7fgeGVJ+rC06cycDaGpLiruUYhJ22o/oP2z
AxX6DRgWcDoYJImFhG6msv28lil129tRlskS3irMnC7t5u9LZNVwfdxq3lRrXH3Q
1XRE0B36LuUeWc/uc/Sv7Jh4BKQPA8d7XeVBV9j9DWZjuEgLhv+T9AoQZEzDCPQm
hAmIn8MxB1vXsx13konDs3x2+9EJf9G+sKwav/wjMs308kmznExvZ5f0eyTXmQm2
IjC8t6ssSSMx65PNZx8hKBMPmJ4WeMkTI55iNl2Xt7Vgop2N4LrquqpwAZatwWCs
vdEE+YXggXZ3Ey5gYpQLTJSKDnjKBUDNg4RAh4DH8vA9/JlJGaxIkIfu7q1joN4Q
fVYb8cgitFarPiGcugmwzyqoiP1yNIQb7HFr2LW6e/uS0edVAldICtx3+0flGOC8
uSVfGxYFLuQ/+BWCCQlDPbwFIU97zooQ1WdcjmzojE9/K7NYPQK3L+v8KVCdW+WM
Xu+T9nuk+sJ5fN6mTY8gWNK848zE/LdZbuS7MNvJGKBVqBxSJLu0bJasPOGfk81D
U9vBo/+/B465Cctk+OKcbxzQTb4pWLKNqDClJrVyLg+y4ChZVx9NtHw9jhaC1rCE
GW7u93PuMI9zHI3GhV7FI6A3sk/5sQG02CiWPdAC5BB2NgvMieu8PouHWhh/Ptm0
FsJzmo/YZX4EfjamCHWIBtu60uBicVbLxXZ2pHjyetxQxrtHNajVymYHAB58XP/Z
hZzsv9n0Jk0vVsAGE5P4wPlhMzn9AL5qIXpKSlgeEvI+8JF1xme06toFsKhViDnn
IXa9xOg8b2nxNtqSepnoUunDJ4uOq13QRDUA6pbDdvt4EoYwqT8fyl3u9z/RcDZ2
kQdiHAZH8PtXMHfCMO+34DeSgjMBoYiFkn5ExOHh33+/60wIldlGTJ/jYQ2aHptW
Tl8BYI1ZK2KsuOesp4AlsBuJE2NEX2R4Yhc09h+6oHNlsQDDavugftC+Aeeir7DO
`pragma protect end_protected
