`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mqEHxLoFTV7GSX5c2lODVB0a/2wwN2y0h4jgCUXg6GoSA3VLd5QUE/eM1dMNKL1l
YO2w7D8q7uVCW8LIgGlzpuDc5VCdpZvSkEMZcGOUt7M4Y4rkPCS4KrAer+YsjKhP
3cjRA+MBBaZAVFYSrqNsrxdPvnI7NU7W+u+EJH0xT+4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2464)
mf1ueUYSizFQsZkkon7Z0Gee+7lmkey7h2v/ReBsU1x241MeqIFOu7fkatm+m7Vj
wiBEgMwMi306+WlWlFHb+KlgRyGk+EVrErr+qWt0qO64o0e+eUyd8RAhFzIktcqH
udb30quvkT//s2N4CagYSBZBQNXbgCogjrK90Tv1urUjmWSpTsf1UL21xzxjzomU
JWuJzCGiC54slx3SslgacSURDxkW1LY7JNvoz88bAIU/OBFlwsjdUmpyyr04H92K
mq6lhpes7TFC5X+sYyLsA0JJOLsgSxlh+UNsRRfc8tvSmNriNLcXgaE0hkB7IX2S
MPPeK0Ug9HmYumfpXjIEEbfRQb9iHPjmG6/c3ahp02Qf2yxjnvN4XHxmZJQnK9eV
1gfG2LZv/OsW7VlHHu7RGti4wr2xyCJNaZO4aRXdYLorf4oXfK4vZ7vUAd+pzfIF
/VzI59MsWvgO0qQR3Kc9GEBUcsHQMUk/VYXi0QqX152CeR2N8rKBC+lbhK4MURGZ
F6IbKFYDYe1g753xoNLAjQpAOrQliIjQeZ+amMD6aauZKPtOPhiWlas6Ibnuqije
GokvL7XWCZXVGTjh29gj3pSy3jotfRmHoh7ahvc7wl4yHNE7kedE/uq96A5jqvaL
EFcuOee/aul2jLnONG3C84j/1liP1bzdpFdSc+uu3gh6RkwHPiHIXUi7S9I8bs+O
LhU8izQ5nam/BkpxrFS+YJIIq9IZsn+ylDqrRkexwnk/sVHObszO7kw8qnrblyzL
LGl6Ye3dvypppcCOQLMzhw2KHKYKITjtEHZypX5CGWqiawrQOUZDoCXxljO0n/at
OFKn/nuFNz6GJmOCHI2LClnebP+3TJMDKHCWbSDrEdlr2hdWCnZkxWLyRDqO7xAc
D/PhsWL7HjJw3kS03ASPyy/MqlPJtar49FyONdDRChdvJzEtGgvOI2poDi0PB3Ls
o3fUilcMkZjSstaU4IS7iJJaXU3qCXGWMjCywGUGxyLoIkhsZK5TW6CO2aOmscYV
kprr0SfWVxIHaO8Maf+oguObyRacWmjk0jgKLfMkSV4OFSY0K3O+lCvMpeL/4eg7
HYPo76qKiJJ1lQrVAfYEkjPZOI14mwcXi4gVptV4LirYoH7l9cj20ImUqQ5uHP2I
NlSvDvR4pCI6Jd67NhNBCPdivcceJoXCPi0bnzSGa/gB8rYxcmt9m7eg7TGsFYBI
1ob2LRePEY2VshyDdCtBXBPsicvoT12n2OCRVJBOgOzddGseaMLEVVw2IuhhLj68
jHijMKKy/LbrecWZuC5MHoT8JCJ7DlAQWgLVSFERIQFPWMSSHbWNwK9iL3bmOmcL
MBgQyDGgeZue41cBLmzRBDWcbAXp9YqihjJbNCELhJGGOhf5/a/rPsd1su1Jf2/h
USwamdx0GR938xKvwl3Qx+KkBy/EKbSHfNHVKeagXzoCLfMA6rV9Q44ST7Z71krZ
b1aZZ9JnSnRxKLr9fTdeE7rukvz/3nnfmo05BBY9m/ibJOwZ5uGRVFLUpSIr5GsL
hhP7FvgV+jEJjnSp8OWihsjj+M8e43A2uiH8D4AqU5KkJrUVX7/1gcDWYZubspWi
VXlQTl0eVuUrvxdyjsJ4VyvR3nvmjhVbOEC3IUls7iy0z2caI2SMAzicr6pe2y3z
yKvJYCenQxNcvzU00s15LhEFz/3SAMPZzmfbuV66li8v5+U5sZ7HLqiiAm20g2PY
nm9ZEEhWGyc1X9IoEE8ucXHP4aJLy30E+e7h7FDC6/uMoeMAQ5ElKDfqXEFhdtBj
EFy+f87gQ/rlbF5dMpy5vTvL1cbhYJQwR/bYEKHQldZ2wojdfejolmZ16J3bvqyX
wHdaygjPyBUVwO2yCfB2smjs4pHMvEYWhNtIjesmEa36Q9ystRWM3c3WU0rpHw7N
dkZZ5EdMlUvGpzLldeADkNjupjEZW3rHqMbrJGPAgVeYhfEctfsOhfDodmmQtQp6
nbnFP0g1Sla7ie6b8A6ngkt2IwMHq7JlF9rqfjbBKEIdiLIc61j33czwFX6sS2dv
T866JXFU+Ds+3fsjLj/CVpv80FIdqk0mjANaCzbC3VPsFx1nRPpvQl810thoHr6a
TVyLsR66rJOj07WZv+9ublrETte8KMQa8bZzj7GmvGKxQWKhItB2WSwc7vQm6SsJ
rHfVVN1bc/z1RVtDOSh10bQEE1N/KWukR/dGWfZXNTr4zLVBTn8k4gbILy0RlEyb
aYaD68notQNJ8VZehsIEPSJLOHD2zQg41+/llZBtDNONWa+OVkDzEAGkFzUsL9r9
4LD6UeOjfWEM1GMK4AF/2jEj1vPUOzKzJe/886u/gInyx/BwanHKrgAGEI2SngFn
peCcBecN6PHxu/PxXZo+VnA/zvxLAL9iRt8ySOsVuVRfbkz5zGWK0SiUIbgs2vQm
XF3e1PHTEhWucoc0MrjgM9hHNPGqWvTKp86BaOxhfUFcSTI8eXMbhzEKlYngck3R
7Tb1HSfU9zQ3DPd6sCIMIRjQ/k1E/4Mf9ZYmU5wV2sIxp3j9jEStLZECtq2I8KQu
RaKvJw56xPTBslOaI7WpVS9DdR8VwldOGzJ0S+cWQ4AZuoB2exh9lbggBBkzcl4n
j5bP9Z3vklp7sjYULphY7s4Qyc1TDaaW4YY6EeYnu6rHvK65Q74O6/Bcdiqo7Aip
zpjH4w0oTlLnfxhejy3K+K4X+wgiF0knCu/wJkyWq6LZIePcBPKvDyl6DTbpZvbM
qqZHK+qIDlRoDJVBcV93U22KHGc5Nkm6q+xPy1Xo5fH1X7twXkqSo967Rl8FbWdY
yoNJGc06DWUBPUz2gbjQSyTtDdk4DnfYoTvmzJIOeOjxgKjQOxYpmROliJZi4iWg
ZVhS3KyvOMuWtzPX46TCkWCir08tzsvXoJ1fikA+kAdLtYv2dgchFxroUQT/N4Zi
C53KN3Hk3x90gz1z4pbfElhU2SuHSEJT4nfTz8k37TP02MCg1/r67tcfpdVaFiYP
fSHVtwFVbrU1y+j/CemN/SVuvPGwN8FmojJmiMHyJY3Us9CtK3M8e9UWBm18sNS7
aogupXl63LOIPJhVqgIeqedaic/KM+fMABOxOoiGct9dJXP5Ewt+JhTxmxSwCRF3
A9wlxl4a08umgon73d8bgOPXjz3eUDTj8VoIgDKF2Pm6gr1Y9OREWFK7qnKT9+Ec
H8S+T5QpMqadbZSMdiu+/iYoe34TdNdFvBhISU6WMIlJmdGOhoneY3qaldbG+kWn
gtaEW3GcrpsRDsh4lLDpew==
`pragma protect end_protected
