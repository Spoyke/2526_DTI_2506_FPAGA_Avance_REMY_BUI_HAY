// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
nLX9dRPXsxviLuR/6GjXNvzOCxwt7VIAFYVbH7JGliRhjR+sAz7sWGq0eZMwh1yJSCPGP9dfHNPZ
AZw8kLDdUIumNhqi+iATQF7xyxZQXL/R68SGt274hLg2tubeRAFEEqnkEoyXm66Ma2+ctSwVr7AX
aRO0bCAGtmuVyA9s24M9f0sdzuaA26zubpnjPMpIZaV9ZOKpIvFchPi+ZJdcOWQAOVA4LOXFFNVX
WAuXvFUwzuGdNNWmosA0JZhnXcFx7m3RXP0twDhHltFBOskyvqvCeL6IvH3OpOeXQaUK0/if+0fZ
1I7dhw5rp6c53n8yRIxEdCoCfJUBA9lP0dvviw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2384)
+J5Qd+DhAfHrUyn0c1rYwW3aFPpJHXCVxlJJyXInH26LeUbHZ/rmJLVVBf8sT7micj3zRrMjId7t
O1fs0dKc0HNz9TsE2Q+39XqVOBzTqUyoqRP802/X052AVB1iA2k/t0aixSPzADvOfIXNbyuBk+C1
C2wwbgrpdbo4FuWffSjRo30W8u5pWWAuLodDLpWYtMMzB7VLBKk526pdN+8LPunYQnbNpG4sn2CT
MGVXwHU0yy+HsIHvQRY9GvVcBLuf/xZUmC/JDS+G5LqGMI2PoK0U6FbsxMfNPAHEcJnO/FtoY9NI
oJ11HBRkQSWv+rvF1998ZTrOG7nllUFZmiZ9YGRBdA9pnDFRGU3V3PtxRz+gOdejjcyay2X2CySH
rqEVih5Uzb0NzGFjRBggJPzvM9AWuL9tuOGn2AgqAUumIlasqlkXYpKQCnkjoOcfYwUoPEaTBRyc
CmL6/FSaLVhCnWBMyqX19iqMLh4YygMUFDUMZLI5tMJ2OoED5Z6h406OSEmHItMw/xhSc1TxEo/A
VDjQ4uSnVNW/ch7HrGj+nObVOCVpyjkwElmFHnXA0HQnmof55I9jBB704mLcLosKDIcaTp4F0vj3
+xN9mKd+CuBi6cJU8Q3KqZw1kTAVPP8x4Ftv54PSKmGy9NK0yp7tkuA1b2mx+4Ez9gOhfifYasm6
fTrDzEugbJ/Tp2ZCGTF2DmWhxokf1GmGb3iPQQcrsqfia19OVY38HuWGT/tCDSvI+lyOOYUM4VwC
WO1mZqAHFtcKU39NSAUw97qk5u/vL2JUkG1MhrCOok4rrO1i6cL5oJdOlv5oSELo6jB3175BhVUp
eZzW9RDFfuV3fPftJssVz7ddVv6P86FAaoWTs3PNwk23I+yNHUNq+KoQdytp0xZIDgPADPsD2r7+
h/LhjjIQvyFDxtkQRCwbrFOY6EqgoeUFQlwn3CKqObAqf0bl7KtTgC3/tc+SsbHck2U8rFPDUySS
z9/lZqkM95nq+0y+PdZD5aFzAw06T6WVRSWUcG0sMkHt/4X5F/nXdJt/V9+zOvrVZ+Rk5ZhU/ZAR
Dc7vy4adPRUzp4axQ/Ou5qsirxaSA4s4R3kJ6JjPN3XP+MsCivtu6EQIsC0fwdzbp0FMsrcAdgfl
CKEjEbdhlayuhemb09jL/47ceOHFVPG01y2JK4cTtxdKwzx069qJzXPEInqk0l/hYomPvW4+3V66
t2uCb84hw7hJWGnZ7qYzPGRUDa/eJXDXxsMdWakb3F4P1Ctb2tQbEZ7rU7Zhm4l0i6k0zir1w3GU
yZpCK19ESRFP/dEMnwwQTnmmTQTVM8v3REPqi65mRoXM+jnfaUnSshlb3WHSuhp3SUF3I1y21SpB
yiynscI/+IWx/GZuFCN64ZDfUKURjFJS58V9NQHyby3tqHz3ajhTDwk05FA0/koBwyEyKVkBnOS+
CqOmKW+30M4xpJXmja0Yu69lQrOhbn/JaabntE43mTqOalO8J9GNn1oBYHOWzhoee+bGf7VRCVrP
u8udkwQhTlppvVfuYzpyWc7iuS4oCyDRDmZLDOcBrKUPkeVBGqFnAsTGVPL/2h9Vjamw1kr3RBoI
VAGtk9B738WBdYj+fFRCo53oO101cUfdPB9oIXOTynsrOZepPWAVwTgfm6zYVOxcFErwCDRqoufS
0+wkvH6Vu0EDD0l9K676QB6czpIA2Gzd5UzGplaxaRdT4KtAB1Ws1dqgmTT1BpGJXu20D6mTxzrZ
pTWNl1gMalVZCQmbESZAUrqCYwdUJmxfrVb+g3ybcAT7NFHFJNuHCzK8N+uY/wT4gRlF8iq1c8mK
m2FgaG50A8OemOXwUGfDK/NSIJAcC/wL7W5rZo2g7mds3xnpjrkPFaZ54wOICY/G+SVHh7y3u/0a
hHbLY4y36TIaZE+NAzWy3NVK9qfFfNnyj9mzFoSSb+yeBvC2YdkSgWqXUrVXAksIG3n8kskFtUhJ
vbqlEO/uSw1I95dh/UDMnVDpItrKkSGCitD8KqsJ651gdyTRrR+NJHSJ8wZmtj1FW9s1iFqhyMHQ
EZCioUXNycyfC+KlPtO/Qk28RZL0qfbwrIzfQQ4+Eg4tE0y6YD5VmgNwc17oDxjd+4iimzuy5vJC
WqgQNPEOnf4UIOXpFLpgwvVruaGxRyzZ2mmsbjVscclW61eIAUQK/CfjNTK41YtfgF4b13e3aDMJ
UASrmMpA/rfl7mAo5q89PJz7DtuKUOLLmSz2MdL/ytAVGxxgusR9yAEUnuGZ1dz1q4WwkY8S/3Ub
uAN/g7Cs0Xi2/9yFhThIl3tzHrK1CQ9kHJjstWPy2qEyJAh+WoXfcb3d2Yu1zwpAOfaJBBsk+SLx
naX+TiU4bK1hJw2NS224NalNutyk2RMSd8en9QBtJwrIBMvOc+53vVPUOYFJX2L/A46Bxyqq6fhv
y+n8DvFsfGcLMCr1qQUEDjr3NqAb8vruqG5aSSTK64ZmGfj0hGlqeOw3LnUl4EHhdjA4PyIQOj4m
uNfSdMyeJ367aphznfudb3ilOAhOJrMw2mMjmqFCZIiSu6O8gFJ5bloeR9xUUaTUMTseOUxcEVnb
2ZQo2MZVfQwuShwRbsenuYwlXy3DNTbh91Jo/vUvlM6NaWA65hBSOMHoKedhEg5cHywTBhQ7LCmK
fgjdJDGRNTo386sDghJT3e2oQnqWAJeBnRQF5G68Ew1umpAAu2BSx+qRuPghx52F4FFu1fRKpF+z
Myc2FsamEyHvoIHA7SZ65/GxKL2wV40C0ttCeiB956sJOkQXc7seKxdqwWOoZAF1IhoWlXNiL8Xf
0WZn9k+MUwHIu+85dVuXJvYE9BmC99ZcnZKxK4isL9dBMFZzyBT4TwSFg5kHRN0mv+sDgvQvW5HA
/pMYx8HXmghyTiX6z/rzLv2DtmtHN69g6pcNkPwPAJiGxIrxRpM0YqBF4ZzjB3Za5yj5ZFs55xst
G1xfqQM6Kd2v2f2banlF1zpka8liH1Ict08a6XTE2E5fpzCXsXI+w5YXhL1e2s44kdK4tmlLJnrt
/SvUtVxNiekXPgyofBoB7FpU4twg64FvOai9T+JRUYQUm/6iIMsDOqwrn/aLu6RqWZ/tYmgSc0qD
Jt2ypm6sQLYE8SNlzAL8qQjnEbgKXJNcfKY2jt6+ZEtMfqx/idO3L4PtK6Vldrw=
`pragma protect end_protected
