// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
BjKxQMX6ouLmZzI3QRvn8UWgUPYTSpyCNd6r8YqLVhWzpqw40dt18AAGJqMdoSWkPo1fJdL8XVbw
MVwE/2uEgmcwLksWZVytHwBFCa9dLMBwOCc2qVIwZddbKRRohoKyb2eFkZzQ72ar6f2u/2UMbBuq
HvheGo2+bEC2Y9kLWUkfefUuFmrTuN+o++omTv/+Tzz7CLD6TxYN/EzqBVT4S9vQYc95q3v0pFxy
rlw7AY4kNi8RZzUMwal8jMUdedW9aRMFGAt+MdCD9yc8rbpVxtQTuVGNXBOsusC6nY7r+ksEDT7V
/eQRh/KF2o05+vNBrL2Yi8m1PLnsYLsTiVUtxQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7216)
/QW+u5h1eyBFBwhe6KMPzcvNvwUqJiEK/vWOIKm6jS0WFHQEzxj/WJjewhqVvrHgDi7yZUBnl2QW
b/jMAYZ2yzkpD5bLfOHFDAmqszFD8wKI0dSA3BnRc1gVKYRHN5QPIROZSv62YxntEwRUjapn6K9K
dCrneLYCBElC1yvzhmD7gAPVynpNnIKg+p81IBzG8yHaUHj1EQzCdo/UgkeJvv66Wtzmvl3tdpOS
B1HJXHlS/PMAHWuZCQ5dmrGxXNvRefM3dPlh2KdkBvPvuthP5faAth53fiAe7uSFGoK6AfcCCnu9
/DJ9I9q6y9xgXH4VIUPJCKsMTlotr6J/SD/LU7IQGCk8ZFQ0fhoAyG2CNsDNsezOZOO5mSi3hYHR
6cY7OLOtLjPaGkPMEh+K8861yiAgODo1JbcSUrt02Fyv3NxFiU241SnM3CAt2z367yvAt+31GxW2
J90ZL1bUnHn7Lf5fXOG+ry4FSRgTQs/ZVphmarxfaz6Lk9z5/8P5K+aWPiSOlCkvX+Uxl3+boPsj
Imiea4cyI20T2j7gzWQ/Tw8y3XXZFMn5sNMg0cZaUmbyRJBsYi2aJKzx72ZPzS7aoLnFBs9V6Fpm
EpmjfK4kYZhaAzYYRim9+L1L344m8EvrNlRivUsuX7bKBlOFYMV5wskZkrZ5T/Hlx0qQHi4YvTww
mR1/pKb7YCdeFH2E/V55jdOIXHzWwPsTjOBaY1NNcXmx/Av3sotkFhRhA/QCfOs34uibpjmK1/ix
Nik4NuoVNbuhPz5yYl6xApFYJ6qiG8t14zICMCKHXXMSIQXcS1zaCbppaKc8dIKqrbmZe/jujp5X
CcVhL5Q7qWtZ3ZXukLvlq/1Y8wLdQim/oNvYtn+GqpmevtfYN/MoDPRyNzezXiL0ryyAWAp7Lwn/
K68i93TmJeZ0ukQeQfFl+bjWtZ/pBJ91YPrfAcYZzB5LfhbtaaR9IllEPMPV9fKfLhE8OqIniJa0
giKZ0NrvGFrZ8lqCZbqxfTNAKuEQq2JiZmen8cM4m+TAc+tj7f/opC8yivwcy8WZBJSnaH2OrNQA
btlsN8NLraRm2aIBlEJ7EnlveIi0OHXAlGxtJvvB4lG9aHq69qJ7/Ii/8+zvD8KqJlBFGBZy4tTT
ADuS9devINMYRfXN1zRTOjA5Kq1si1ShNULd3CYbajlHnYq+Bdbs1OTjnzHRHqLT0o39OkrYWL+C
mTAAMApn8tn5jHzSzjcWe8ayxyCJNhCh1mg/Oeq5EP66+hEdBnu2WMN6tJSe1nyeYRMCbPApKLc6
89BHvTa+6W5DmsYMgQ4DhCRWVD+GDvgiYGZ91GRAJ7MsgQgG41kvoWOcd66UMrupUfi/q+KTHlUe
7eSraCidZEtnMvqtOgEAfBcJMzeUgcb6WjDkluxVdUWDlSckfdvTk78sD5qck/OoiKRKyovs5+RS
ETePcqH1EEU8MMEnxkJWgPBuFDtXzNFkMKnvMZ+eW1W9o6sZh9hDt+xwyg4DFBWLdUa+mdZfJg7k
+KDBLN5z1pulXW8HKZOdngugXW9xBwuBI9zR9KU6RdstjaigcAURf1oQ9iDbIYsTQ+7NNHLFeT2r
CRc60ELSVF6bOgPAQsjqN05lHnLrb93jDgHveNBml4ftSw7x5TIWOCCx/S9vEZQkBf2D90+tu2tW
YadSb25enTKI3QBQ/98C2/qS9qQH1GLk+qJAxEcl4NJZc7kx/wUWeZjctMgUG1+C/mUNMLfcu9LI
ulfGaVlNN5RVEJQ3dNPPbH4+ThoJwPotNYqbOGp3TxbZlZbesAUaE4JmgDsAdFD3Md8j576wohnM
Ho1tfoJ4fIacqok/WKJ9mADmT+I1uBSbFna5AHKsAEWdOGrnsRof4FIG8yONeh/9n/LER0KFvlFY
9qUApwjAlcEbrJwFqU/U2PK8MADLDGNdUKzfVt6hpTHjPOqrFSYnBMWSPfm+mhDibLrM3tuxx3rO
NFYaHJamDl/L6Zd+nZD+9VlnzF4cKKckv1Fc1qlhss9Ad5aGl/qTqIZqeuYGFGWOwAb/vRH3Cefi
irx3pTVTMiy/i8V0JxwCuXyCJwczS5iYpIzhs+9dqe68/3d37N4U6ZQnYeZ7g1x0aHXQgkeir0t7
F9c2EChFfuBcCMCvsbrtQkft4YHgAkZo6xO+kjIRVLWX/E7CrshqUtKEsFGNjP3TX2LayCzYlAiF
ND7XVhG/Nml1GhR0hsr8q6qSBbVTJVnxtYn06rKavmX1CGMX7BtJeXDCtQToDVxpiAGyUAYNmM6S
qoSZliCjhMkH0GWOI3vzmUrb8WD6kxG0uOyVTRWPjmF1kOHwA74fNgNGrihXayK08Kq/XuSurvjJ
vLz54cNHnLoSk5XgKHZemxQlM5fEtTE0QNsDJJYpegAPdvVqwS2Os80atnLnrD2irdj+O8wQjmhf
WwHNmLdSqELQsNwdqrJVpFopEc+7YRO5rB7MUOeB2OJ2fLdW3yh8qWVRHXXP3bZxhRi4KcCn+Pkv
rkE5NUntzs5viHMHsc0dzL2QKbHE02fr5YJxUy1/Z4W77RB4GJrT7gmrcVut8CqyZa+R1qSaBnyo
+MJrVCJV/MJ0zf1sHrHhVee92BrDeh/r1ziA2Xxnbtfk6F8joYbezISLCkqn/g3k3SEY5pQuI5TQ
asf8xwHksFCPXxFnKQexRJKVxvlGTqqDm1KcPH5HhxzZ1BZ7jBP+7AcGxQY/ujGUNV+hpKFzf4eQ
ahf3EWZLoZQHR/7rUD61wqG/cuNrMENpXwinkw6zNmLRCGc/dIKqoa136uOHLwJzygzwxoafhIO0
/s0rSS1kEtPfLAynDFn9PR7xBnsnk+W9BoPRmyrrVrgaH/7u4k2jh85AJ7C993DPkInYIPK6Wrl3
8EGSn8EtxnnpEK0dL8wxpBDn9Cni6QtWMubEgzSNWwGkGUIaZ0+dn6EMks6IqyBkp+fpWZp0LY4X
5xamuUtV/5AdZen37IgSdHsxVWEeF54XKSINi+wt993dKn44Ta3hYKap1jOZTHbXvmFoF6KJJg75
tFTj5kpk75RbISwXHr566CYWzYikMiqzoffEYKSexoJeldyzeIzjlG8eP8O4VC3z5EgHP6/dsDub
PfnwvVH9pVmylf0nuuKrET/9lxIfAqS3iCh+9NbcN9xnXItrZhL9I3MIirI5lw2+6mMDopHv2bnY
xiRVmg6hRhXckpZB6xNSyPBtRBHY4CH/wLYTt4iFEGf/Xdz9HnEOUKoF6V1K2Hf+9nhGyEmbkErI
xPlzQFs15hbq2dRNE0KssPvblUJ2B6o7C9iCDIMSAB8+mTeH/ItBsIybqzN7uyDGPumyFuX+x+4t
hdNYfDMPwr0Uza/FvlHmWgJSJc5h/HJkzN4qTYMAbcS9FWjlV8lmRzb3CDsWQcyAA14nd9JM379M
pShzh7sxK9OBtG9UVVMb2Qio17cgASoWLMBW3N8OszKGevbZlMxzqcjHi4UY9k7BJxeccD0uKmJL
7kRvzUYhu89zuwlFNKwBAsDGoyBbVLZj4VHYAaXPAKzdqvh39z31ra2c3N2GPMpFVt08X7VgoFa5
xY2FW3BdEiX5qYPAO/ZOK/3f3PLfiTwaPnrBzRTAkrZYabnFwibGnpxHOgB2dGeDstQ+EXcqVqQy
fhgPfF/xIyc4a8uW5e2vvwYSzO8ZCkLtcougWLVORhNzO5qDAdhNtzkXixxV1MJ8CVdChYWlg31W
Y/9W77KzAIGLD7b94DKTy+fx9L9YM3mvu/fHnuXJfkBrVdPavWd4NaUPsV+JrXbZXv7VBkdqTi3J
FCZpsxh37GPxnYhjzbDfJCUEvPYYl04UMFidvim8M89CsejNTydgNd0JhvXlzxObpH8czd6FAvqz
iZVnzReLupWBWqZoCuhN5g5DcIAAkD+Kam/MNo96fHVqzURVwDmdN96WpS3FLQrtzQ+c69Y7/Ams
l5Ua+epd1Ht0/me+0oi8m9S/cbaD9wzizrLS8uMg699CEXW5YyvMZ/vtDgN1GKkIuusNVjqeeh+e
ZyZVJLFpjq5q/RsKgMn0NetlE1XKgWSyXPliRjP126oIcNka9lMhhYT31R+k4mnyJAMt/Fn0a6e7
wzgbZGLcSDXhJPVVL5bsYttXW2GxVGd/S9NOaQP1WQJErvfV87WdWbXbRsP41Qst0Zwd8cyowIMV
qXm5XzEzJGuFmz9v/5PlYLRvrfxmL+IAqILSquvdkGNav6jq8xHDKoztg7ikd1Be4hcMaivICLhl
JkOhWChevNRCWx5l3VzbjFcgKeFEtgxDTeYxpNbWrdHsb5DE5OP5lp7TJ/A1NvzwVmaGd2nbRY/e
4aR+xc8Y9aU5jZtOHFwT+HjVPGLFIQkr6i9iYOcqDDDk23D09AE6UcZpwb9oUzfZuUWHdeH8tmy2
olK7l8GewocbDLpmx3Mh3ffEB/HfNuxxHn87UKTA+nK3iWFflgdBunWTKi20Jh+IEkPjdUI8DuDr
BtHhu8nvzqnHnTnxRkB70ZMMFkBw0p8L5RLNp9K3Hxmnnpv2jVZQ5AB2Uurpzz78Po7GrNMf+ULO
tSoH0vRDq5QdQD+ZKvjGSk3+JEzxbPZ1P4BkfHXnDLBEHTYi5qitbmMFAgiOXcIpg0ugMD+TekYa
fEbtdcYg29Vu5sZgYxNCn7obCl7M9eT9vmr6wXENt0dUlZZ9jfRIGg//i+9X9hOsbNyV57lppeC6
BUTttzg7NXxLbqI5AwQ5jj5oa8uBAp3ho4y+AFgBMT6WLuhjAHP8yOy34iSrWDnWPGNM5oE/9qOz
VOlexb6YT2ACXKGrJXwnmizHl7Sw5TvMY99kqEKizdxf7SfY5dZ+f7i/O0rCW/uWBBjI6D/VQJWR
5W1nVhk4oTpWM6UvtTTh3KQWg3DS+N2Js3LNgvKo5smnvXfpFzQUrnr3lCvJMFx/hkXpoOCf7IW4
J+guOnZi1Om/b+9kVx4tI2HcnfvFQkGLO4ODUgX0f/W+38Dg3SHPHRbITWqiDy8xMOJgpo5vqS4R
ILuwne4tnxSrTqviOI8qk3XSAqMItf6N5iuOg+L72jPOaET12/HEOnZ4j6/8xAilIzKqbLrGe9Pb
L6WHjUIbpbeo4ouo5rHLy4uBu6F6Ort6EU48Rnlqkzu+yWzaBymxCsRzPbCiQ8M3npO0yuFOF1hl
N6qhzGwuapr9qSFuIR4TdsYlKVnDhIPdkc7DyFqLuKWC32XsDJQgRhfbsvSiEnWhLFcv+3k62w+Y
hvuWhKL/J5O+a3R4yyNkiAKy2qJXlhpdAxUIshiZm3P9+hEH79HYV0CN/k22DWGp+lCeTasnEqCo
fmHE4BGW8z5f3ggOke01FFv+DiexDXX3MXno99JDSJ3Mb9s6FNgbGLEX0XUGgz343GzouFY3+lVa
H6+ZtA2PvacMI7ptlQQrlj4hQUM6cad3/QkblenCkAGZhImI4SCMHLLOrmkpo2kHIxzjLnLoJC+c
Pk+48mbvkzphMpDxm/DIPBfMdUHV1VyYC820C6cl6dXwG40SrWZeiWOKgT4UZY1pSWmdI0PKCewE
P9Q3qJqd5zKQbtxe6sreeYjITQ+FzSM/KrNfOLEYxC8mGZ7runfsHrekMqANA4SdaFn3tpGbSEKl
8xASwxpcBFtkcaITMUKN2CWqqR4pCiiFpma7IIKhH5j3UE6dgQi0BGpTqp5FjCLNHuku2rxR/qMc
uZz8KAm15rPkV/QnFqF+ZGOSfDXMHhQrCoBgoxGbRbgxz6KZ/5pWuO5LWUMqbeiYPYVcWFFxHn5+
NZwYYPYFGDL25Nr049dz6gmbnknMFfyQl9GpO5v/sEKwqWWSBpD/KawIQp20R3iaebB4tydW/bXI
LdNvqIAmldU26R3on71C/CWWkUJRdp5jy4HHj/V7C/705ezXktBBqug5DGLTjxbiBA0gcVmJBQLt
pu+RvI9whqkx9txruumfi0lsN2ztvRhrGhm2ZMDhslPctfXPENTwlPdWrq/JUgqsFN73LDx9j+Bg
aV9cWl69CBD54OuHB3yzuotQ26QlfygesUZWsS5MJBdT6wKYKe2b5iqspH+KikpqljbzgQjfBH5F
jU+Ue2NKOR3uSZphFizk/hvhLEkGZbwiATHiOx4PJvObYDK0aisUXzOsWl8n7ImSCFtAghqExCRx
LYo0r4FCyqp2oj3yjrQiDSZHFJq/xA+X2BnNw1R5ml2NoWytQ/r0zDqk0CXQw6Cx69W+ICkhk8jg
qgr+Qvf2n+s7+f3aO7kqNttHJ8+H4kQleaMio/szjEcg4EqtAyYvHUlTroiafaJC+g2vKTuMzq0y
o7WV92+hCa7hoilXM20+7xUKI5gp9fvvs4Ynn58xK/oijTd8/LnbzMDF2qC/O4I/b4k34F76n1HU
z1xjeHYdz8llKvDoHphT2VwG7d7cjfxcwiDY7/vNBFgQu96i8LMgRnpOtgMYTdzGMzeTItmybQ95
x+AdVdAnHCKh7xUBZ/sRCN2T/D0wzHjZ+zBdioUQmHUdvTnwJumCWuHy0BKnyuNh10Kk643aENzj
v7hdaKrj6QNR23MFEV67u+eyEvyg8EbLlXl2tWINndVRdd4pa7JWXIAyPjV5XmtBfW1h90xNtGxX
qBKBc5/FxEH/oAFyIbWCFfdAeT3IqUb8fxfhXSHqGpzlzy83VdbWRDGcio/dKD1pQ7r4DOaJyC57
+qs5zdBdSYQlMNWDH2kWTwql8BS3QiddfNfXh9c21ja4XhCeBvjFtl/STf4c9DUzsnil+a9n0Jgv
UUp8M3oJmoOxbz6Ut//LkL3c62dqvkmXhI85PHn50yeTcYQAG7C7xCnPTEGHiEfosMD6voEULr1c
AK8/wS7NTuO8z8yLRstR6K0/dc6PHu4o2zAHfJGlNj8XAIG9phzZ+YSz9KmhkBLr9U1r8VVEbk7w
SQmWXbXHt00oCo+9CJXflBuN5QLRxbHFNYQbBLXpHoIuQzOX8qZqUdLAbvd1CD4sTYHePBoR4l3w
5bEXdsq9mZrcLZrIRFS2sn8DVF0CIEX2cbyQ2ODIeQQnBkB01N9lsqZYheVvkaxynm9n/RkSFS8Y
/x6oL5ieOhLfuH+2NTKQk+ImS8Liki/H1QJPnilhGvy9rmbC0ysgqW3QZ3FLV301KxM2iyYwXGKo
QjjDspzd3WK95Bj1bpcmgjxsIjGRe/vFkXClOwPxrQwwieWihPwWScLM73synUuefQBKRKST66xV
0ewBiMXBlz4BYTzg3K5Q0wjmroznOTr38is3SQG9a1yCugDnQwv5o1wr/rAtYNY+qqn4mUnigVmb
Ke2ypbE3OkjjymrsNzENNl2Flt63LM3pgXimy2EbgKsptFNQMkOb7l1MRsCboFK793iOOKaLs0cJ
nnb6YTP96THBT6Prcoi3SKwBF3Rqj8WRSpNZkBHTG/USMkIPgMfgZ/FQeN66+ZvFfeJRPADhcDhQ
4zUt+WlKCusYLrQKMHDtC0uEZnb8+UQlNMzhhqllStNB1uNRU3S/tpfVDPl0y/5ViEkRgGqwRiXp
P1SB7LvCbgq5Hp1bbVgExItwDTYm1DrDwIKHOEjM/mXrZqDJondp8OZ1sWPIPzC6UwWjsLD7xJGO
MsVNaNrOYRsZWf5zisRnw6/aHEx43nBR0RgM4oZOhlcCWBGUyg0aPROdxnakJuph12qNjB+lAG0S
4kMN6PVuNgO9jUbWFa3eA4zziV+52Gj/yaZ5fL1AE4NKtpMAibxN4avylKdXSCKeaoKUdh4wpKob
B46KUWi7Hedp+l+EnMD/NIWuaPlCPxQm35oHH8WC/X4grAuRcS6f88Qspk4G/VJc54afRd14KEIo
bmnhJYeLSgZq9RBSI7CoxXqbOdkMnFhbXH4w8n9Alm4zWTDje1W4POS+Vn0Mg0qu1D3FHwp8jDiT
glmi1a5j+9ftsDBncremYuV76REyvJtHaDxnmpplCGVV3fEEBeAGUo2dVeh/X1uTb4FiIGnrINJi
068d03ifxY70+maYKJUO5oHzAYMFR174nacx7D+f+HTi9/0TJgYa4jGv6Zg0yqa299C61OZ66oOF
95eJIevf7UVc5pHJ+ZvhstCbHu7UbO47sIwvohL5a4eYeAJyxNj80Mzt2PWrvhxQ9q8JFHmesCzZ
YRMR4vMkgYenQKVUKh2vM04eqhzUVnDur8NXBt/1M4+yu92vcxbr9E6q1wAXbNG1V9PAI0qN3JVW
sACPcfW1uWJOhrrw8wjkvYK6XbSFcxsI16ya33ZwnIDv9w6s2HxGnDecSrCfv/H+C7vBBGcUFPd9
yvwQsaMrMem75EUdRQsXZRJncTxtmD9SGlRisciyZz4KpBIpr50CT4CZzH7seD+I1oEaChe8At5Z
JCaIXE8aIU+OY+aQsh9uWmQ0qZdO4GwGOGoOvH11yAMVR58/52fU1JzBRJqk96+TG5gVL5NhSgUe
9uAKlYxUmKwqq5Af/JNTmqC3cVD+n4hzlQsqZ2vmRJZnmwLHwP75t7tyvhabgV+jkAK7VLuAMCG7
rBFgn5QG9vuj1+3XIaqc+wLgjOH83nifYHqAtH6NO23uA8xZ0HJcU+WT27KR4ix9+4BSwmekM/v1
8uPS8/Zow1LVXjhZNTYryXnZIaRfQA8qqJG4TpgLoShLXVFP5K13NYM1nuiirfjKSvHBFgKC3J25
b+w+IBpDrHXEOCDhdDebTazStXJblvcl0+0Gk4RSZ63/YtWfMNOlpRRuJbhrUnCSPzkgikmayaG+
TTNmLVIG9om97QjC/pca+/IhVqd+3EExOorQyTfbRvyOIJG3EDCjOwwpL65wlS9vn+SB+ws66CTf
mC1W0+CqTSS1NatYCOwRxm/geP6Pqp6eUf4CbumFwymTfcr/wFZdCImvFGh+N6Qt42TI3Qlpdlpw
SBBHPjnN/kLVZSERxe/8OTlqVTwJNM52eu5rU5gUn/PYyQXKuV/CvA+otsoibWDq+8xjdScYGpO4
Y4o0O7LoLMZMSh1z6Z/m6BSFQMpclp1HGawqUaBFXzoEO5t/fOlELR0dMq1Bs3Wkrgx9nhvPNsiX
WWq4nRXtmWlDVzEZWJZl0TdGUOCXNpLwRCoxMktsI+0LhVUG33XzuXNVoZsZvzzaHaoNKeFTz+hk
fBorGQYTAylRmZgBxzAnM4s0gIQvp+tPLY+tZos2ihcHtHePel4XeltyFrg5WSNWVfE81eapx7rM
OAaBy01A5mB25o1hSgLK4nC7MZmcT3Jluix5S52mL1YUpHAXl7xiuYd9kJ6pvxX+t/OK80fkb0IL
qMewY7YA3e3FvclNfyNv/VfbOy0k58Kym4wRKhwkenvfh2K3/6/K3F4W+xdheCjFAXya8rKHgudH
vI33bGw60q4OgW+tLsPoHRlF/HgAMA5b1eLPv+60AGm3t3gHei3/Mt44DK6TiXLm8Mgxnt6RhvLh
YNntTH4FegYmFf+82LyaQXnc+po26UKMKLHCeq8j9FTIfJ4yv22yc98t3pGc5vV4VnjBwGCbKutv
OT/F1gJ3OXOQ9hJbtXYAo5monSbd6DjJ7SdsZz9UR2Kfo7lYFGSrEgwMKjOuazulh/BrwKwbj2h/
ZmGO8pI/fsKhN74feJwpk3+SAi43H1rC6kjZNfPcCa305Q==
`pragma protect end_protected
