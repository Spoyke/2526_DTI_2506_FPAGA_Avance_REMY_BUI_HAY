// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rMiryjxSQh5YS5VPp/0gMN6eGGr9TNGLg3IGxQB6LmGyD6IXgjScQf1ofJcjMCVkFeT6JxcNqVl2
fAq97hYqguD0/YztSPtE6Lr01De42cWY7ImOZ4HDbmkwZ3oz5wTj8Ouf0oiBepTrBuzDeD2YHCi7
/rn8aH6d4AIo5hOSRfpPnQawmr4aTj9GOFNFiLCmOKJFO5PkviPWNnuVH6sRQurwBeTqwZhDaqay
2vt0sgLWFxP9Sv08Ll5cdxkOgKcrK8SpuwO7ETqoAzb0yccD6ZeXtPwXuGaJsmQH/AnZQN71S2B5
vY6B2mH8jRgh/HrBfbVf7/90QKct20i1jJNTlQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8960)
JsLIsznbPei6Z7R02CBIVzfAy6DfSST0GNdjnu46dE4HVLN+e61WloAF3plvIiey3mSzhdIxvBiP
63PQHRbwt5Q6oCzGh2+vP6tCszof9Qxy7o72kP2Fb0RxfKQZUaT7iBFCJf0TbDnSXYtBsUMIe7+M
a+mkn5fdAIRS4vsMckz9DYFNmY6p8SdMix76DhamuhK+QeIqbouECjukZEmkVQc8DNogHAbSHXuI
8T0ro/NZu03dpY5nCREt9WoPsd0IafoNywFd/dzWjZ2LV07nXp+pHr8QRflcgimBdnkZICkW+rd4
INcBlWbm9WEwhdMTG6gqNHu0HzuZhKereP1F8OVgDw42OvFeiJu7thM9wtS3JwVUh6cSH4j/vbpn
PH029YEDUU/gQV2347++3s0Syr2wmCQ7KHyh4EIDtRxYfavlBpnDoUvNmaPxDaOH2xo01EIJsFTt
6GyET51fATS8MC8PADFhQVpZgGJHLUWltrD8641Etkhl7AGXEHKf/LCNXqs38Tq2kXNrbHxr7KsB
eJ43h6VUo4gM0UIE7/mTLSxR21Rh5AdI517ZN+pPgIhX6hRQb8XCzy1J3OADB9QdT9/0l4RdTZ4V
K38oxNw4UmHNXEJoqW/jV5hJs0REnwuW1oZqWRiMj9w+jUBCk+oVOK4tn4EVmH/VYOROHDPgd+Lm
/vJt6fEDwqlD2Vb7EBoJxsUZ6I7vr/tGM/SlGmaj2GCCYzJH0XbDw3Ne2Cyj0YysHV7+fPAlPa5r
jCJhpYeBwt7cRsafBST4zHxFRJ04jAEgfQJzEnRI7Zyij1QmwNr1K5JdxsMqrx06Cg4VfHqTmdqE
WFctIbQE+La1DAQn8QaWkECwFOob9oszZF9q4CJ6ytAEWRMQ682Kq8XwfT61LMzRtq4NgW84JJBi
cbLFTUTjaBUE8jh9NYOURfpXOz3ZqbteXEDH0MBMxFeXLFYpFWzrVhyY1lEQyCukGxpQce0oRqkA
XvM5Uo2mjImIREyFKArnIK7lYp6WppfTdjw58gAxi37oYx9aW9wknqy0ZXR8IYMuL0EGsbCTAawm
I1tnz4kH6U3ThNwi3VUoutyv0PeJA7yu0jSSsWkUeGH61IS7OY2unjzxIEz1dl6ChOG8GSDp2k8q
x+qDAyUjXcW/S0+SmpONbQsxctR7KzD493CB5qrA4ASRdiuhD0EVvB5WTQZQQ9ZATJdkiqwmU4oq
tLtbndVyWdmuOqn5W4JnXkp++JcLCYWwmn5RpmGvjUQnpyuEhOytMF/kdDlUnGxIiaXmgHHXA8Hy
Eet02yqAnu/8a/XK2V0Ipun0p5VdsHcUaKuCkGO5UyBIzpzqt4a6FngiA432UrL//38YqnJmRx/I
aM0tNfuZvDsHFfhOX2KDDFRnyq8o9TypMvQTq40+3GKF9vjDPuHCM3x2w35GMoaOEOOBReLJUjX/
8yRxjA/08uzyeaj2+jkcpFDt+EDabQRkh98dDeFo7dId7pSnHdWFViJBMnLc832Kc0/n2Pu3Qz+p
1Wh7fXLQmO64kQpjsTXj81zTelvwjag4tKn9/a9jI73T1I+3V8a+OtkMRjPBsyoRrKEaLYeW6DVB
iWeOpAiXYQV73dw4VQH9fzOM9yFAMFysteX2+2dM29vpKQmvbKVmz1kC//F2hep/jDQWgtihH+yr
bs274wOw6J6iocGqOQqlrwZbpDfxXmE6YkbaXbzh5l+UlWPHWsvxTuZ+JlOujO2sKGqqqw4u6YWm
f/F/p7sr9JmwN8NcU+w+jf4KbowfwKNwfBCjAbzhaX0EGm0FXgsDNj8pbYwI3GOxj31DsHn8Keam
xbNA/yKQKsEAkBv/tzzy8euxqvl7mLaN99Xh5nkfCtBGmIh99LkUxUkLvyIjFe7/26M1HjVXhdoB
WLbvjPbKPjSq49NyNgAIfbBXcABj5nOJ8rhy3Y72cT+YqN/nyaitAqeDclz5lnEZim87QnQgy9qz
ZeL1uhpoUA4+b8POwfkSYWhscpEbfPqve0ZAuIDpugq8X0ASkMOuchlJKSx5z5AuLasVyERXxfFH
WOEd6LAYQg6OQxyoJkfG2Ws0/oWgdPFPsw9lKPm/zLdPRT00JOU1FpMJlyv0I6Wc+NQMCJDkEhts
mS4qC4CqPCWolFPd/uV2BqyAH5kGMhnqLCzD8GQVKxTNVHjCBsRK/C2J2Hy8Sgh+WYLiy7csJjsj
TJHkEI4YWAYcZkFICNiUeNY+D+VcH77LHKsCMA1trVnPScyYyNO023KsgDvvE6w+ZHHYtZyb9I0o
CaaefIWKtvjX/iQZSMAyh4r/Mhsb7FWC5UCi764d1010eOHy2hgNe5YPPKzNxS2bIrHwwDIKQHya
M7IB28Z/QO3f6x+AQ4soR0vAlYUUHy+UwWoOyJ9G8DjfslGX4FNb0p7aAAHRos5HP86FXTp+OE/+
+JUmb9v9G4aGRsmYryzZCXiFkMGTttPMRIgJRklAYjpi6MNFJKZ5iyBMXa6ZpYpwAVPn9G58L1bn
jSkPBmta7RWQDyI+myIrU5Nz++otfVBJZge07DRFmbKStTeEJ1NCVFR94Z2alq3EUPKebTPZToRR
qgwNXFoe3+IYZ5AnO5togP9TWE1GMpr+Iuo31UCXt8OKO9ev/bMz5vxZNX9NkU7ESaRc/h94iwc/
vFVQtV9oFTQEIbIuvvsD1hAXW41iJLSzCr8L271cAU8D8/h7SDs+kobcHFB/8TSi76gkExSETDxF
JF6iaGB22I3tTl0T8y5hKINwsRdDyToMGyf2prwvgQUGkMAjOCGNsDbQFaD3sehKwixHsYG8Lj6g
wQphPwaW+re9wbkAIZ5JcjwdIGCEfQWgbzpMW4t6WIrW/DGSKqcI82bqhI78JhSB+gw3NpnT0DjQ
7MJWCmoWX+M9bDBXTpmeiTGxEK0ACz9C+kWAYbXw3UhIj4U6RowmPMkXu+dAbPam6RnrMtA9HQ5B
QvXdsvSl5BBolXeySNWj3r+XexC1HSxebW1un0vzD6CVhpbcYgYW+fvRigz6FKAPwtsFc1D+I0+9
s5GchI9kCmOYASxDMzg1RSjt9QpT+cKUEl0TE9ARuBA0I/jsHK5bd7w6fZx6FA55u9hKAJhUM63f
Gq2YJd0XSuiym9Sn9uyNZk2NSbH6IqbB7muQhkX0hHH7a7TiGeMMlefB7MeOHfQAwMUw6ZJ66fmG
JBmHQvAkD2L76tJRWozrbhkS07zrAbeu5PbFP7UyJcrQcGEFnDm19s3fMvaMD2rcc8KsIGPhLCyt
xcPki8CPc9/rpb23DgtL/nkpKyDdiNaH0tGksPJRuwv4fEzR6iLT2Z48YAa9Qwot0C9+2lYH++Zq
wmC9m9ZEnCvN/5qu3oXoz9PBiV5UweQ8RJfbedDShpyoGT41aze0vkOOO2VqoqRaUdV7nhMY5RTo
r/Z/fvwI/sqNmaxZIfGr4CIYaHuCwhWW+qkRZQQemMBFsBogFSAxWHJ+A4P+OEu4fn8lsYJiLviR
Pkpgajg2B6pUDjn5/TeAOfo54wnswN29C3zjBEKwJ7U6PT4O52JM1X9OIWxQN1lkZsy9aP4goyTK
OtuVBE6aP+5kEE8daduTV2lJI0iW8fHu0gxEiv5MX3Q+pPgCHGf+k4xLANa8i2eakEMAnpFKSUNe
xZK7fwxT9yt+yJzvgjSrEPniRQDxFmdgdkHRuQuVaDHuetZ84y8N1EsVsumagAXsowlDGfndwe2M
NZiQWAbkEiTH3e/86LUTVfV1soFrMKaHLc+AJ2nkXbcOXHO2iYyP/NjlUlgI68w0hrQi4QxJsKAE
gLRazGMIo89HO8IFDYoG3Rw2tNtFYRv9NUHXoC2B3mMQmXZNH4qo1loAyMM9SSkK+9x8XFaqQCXC
f58XDqNROZgBjis0pObp/BzbgpT3+aFLxrpA9IZBAjMWnFDUfPPRV8AEXeXsnrJqjsARCTpbTv2N
YPtF/DOv/rfJNfkAhw5GiR0mc/obhg8qt8K9RPjRx4qitAlAuQ0q2fJN+6Dh3Hx9erbH8xezg2Z6
3JkL6dC5fG6090hfHxCV3VGxszGRbUy6gMmDNb+kVD53p8yS6iJq6CFUSEDNyYihHcKWJ4OwF5RB
HiefjwGGj+8N4bQtAUNIQkx3URNxBL8TYid35agPLRaVh/PDQ28yfPWgV06ALQjs7OxJtmsAsshl
972vA1u3fAmj85blJJEtBnJTXxDLd/xupp1wKvU2vPogOZuwMMv4TjQ39ojJVlROL6q9/bO7RWe2
u0dXnnMqg3fLt9MbcpzExxjnRsVOf+80PN3BzCS8Rz74G8cMN4SG4CPkm3XuwYbnihFYkyFYJ6Ts
7Ref3YBuBPhJaMxS7uE3pT9xHj39fh7crky7183mVwA/xF3BFnDQckfMZXRSiXzs68JkeeEhNy5s
BBQ2ScW6cxxyzyrf9C7nK/+hdH5n7ai+yheqlA+3p4onkqOahPE9qKfmyr5jILCLPGDkLIsW7qVF
cPo52koExBHUtelkSUxZjud6xWBo9A2ETgrLttyIZd3DQp/8HeenMdymttzR7v/soHJRFxXbeAWs
GWoVput6ytlUA8YjWxuvTI8QcGIK31klzTXxYSH4Oq/MzDni8sPoHBmLvr8CVMIZpasxab6zokv1
CppLnElKgspBvIMqZR/41nhvtj7bKVy3mJDEQSUsYwQElXWfKZaVw+jsQTrvJfvZ6Mu8gZUFNR6l
5XRvVvZWzgsFJK4k9HFRtPgVihnvIZBeocY2IlNID0t0oGT3zLuY0K28zTZgD/Ub82pPladvmox9
ZRAFu3coHNGzUUfF9kc6MyOhZyq8EkeKyoOy09oig8RUMd3AV8Z7rHfrpytuwFb775/V5eercB9Z
tdt/VVKEMMLaiVNRm229Jl5olA5C1pzGTz3lps7SRZXyZUoMd0lyLV62QgXqKXv48MNAGXGxXLdL
Jol2qH1/Dh5tXR8qY2l1khYDIawEOf08ltSbqn1E3wYjLIvPMMmCh8CBTH8Xw2d8hg7SCtrgpdZW
V68aNlIg7fxucOV8SXNoMmqHDJ+qb6EirpcOHD1SSqvmjBjESScexIzwN8kkkCNS2ubmctjdPOk/
cXQ+HDkHWIf8cl6lOA/EtIsx/GdGpFRtiEpLu2zKPj/UZWza+Yp8bLwgCnTwJdHnqw+3OWGxxiqr
glwOFrgoo3v+/4r8rb/gWxe4/Zk6g73ZJo5LDfgkDo2vbqvkY8ZnlJSX+Mh5XTsz8gVPOVrA2LQv
REN7MVsCe7B8zP8OH+kqBe6m8mh3nxsxwqpFMyFXLpuV5WT7UR8to9+t9G1yp3qifkSPHfWcfkvs
yZEB2UaC18qB1HEj58sk8QaL+giAJyYRgOXi1WdcQvO4EaFTppHPky63fl5R0LB/4uoIgYNTSayi
J/hBrP5ajyWbUfgXz4JKl8M6HEZ9Uk5bf8e4M0qDa56tOro6kUn4Sl2630kf3SXhTEMdZVaeucgz
VDadoAQu0DTCZe05FGss8hygTOGam4x0OtgQqZXlHk6yRDkyQZQsx3BSjmNWXDhYZl8ojaxSUDj/
l3wyTORiCUHIQKyStlOl4voLeQEfgM7OqXRCmwkavOQuZcoCRGgOVclAI+zRyKcp4UaAPffRNNzs
uo0e/IdWRnSSAqWzBkjluCmzrOjAZLjzCDGenM2kbsmVwR/qCcrhnqLYLNf9Nhy+ISOIBZk+3cLV
5g0VjCjQtjVNn4gIpj1CMD+6x7S4a3GjyC3XR1jlXN49iiekwgg61GLZaMBINAT6BR5KsYipTxtT
fFstQwnesApkmpnRFuOb3qV8ULkXImJ7ih1ZDgabKKN+WSU8IoegzP3B42ZsivZMhR7RZPNZH2D+
VOD9a0wR8i2S4A8Vnhm2LhLQ6xGlDEY1wBmjMrdnMbidb0VaoyJIt5IbxT2GHHJD/0yJz/tgQ/7Q
JyCthy8Wk1ZzoQeOPDwXst7frdT78bTOhxGDMpEXlwUMmR4wjej+OtLeK74pjdVuUH59H+6qSEmT
1yDDJYtnJXrJOvAKxJOAEBvwkrgb2f6AJH4eaRDD6/6RiM6vrwZChF2HICXIqDBhKd4uhpGS3ScC
XSvJEmDKmUdEIaCTzY7NKBXm8iwt9xr7EOU4NdKx8Y6Uv12Ss3cFd0po9Yx8eBOELxbS6l4V2i1+
1i96xWhEx382Lw0Fwidkmq6m1gmPlDirqrQrlRb0L0pLV/MRtJ2664kG6DJHQlpqMBBCGFtGxkqF
GAOmREcPezVL7fxWe9g34tjzvqrRhEhzWvVkHc3jSFg9JHlEnC6934Aa9G0+cK+vlygfpM32HjYd
2qQta1WzRd5t8s51VB7U4R2Hw40xgrbQ+Nu/2XDzH6vnjOPbRmE0e2hK3UiApuCwCDSRUiT4OCW1
R5Iwc6z8KyitZDo9Z636UIsUki+kQSSq5VL9J3CqAo8nnn32w8EQxElGxsyM8BF5bnIaA6X8xRYM
rQzpN5YOgcOFfIg94ARIMxYkRJIers9uR8aj8IXgDpjnD5eHcSSu4bC6xXojo1xtrdcgmjl1TvVk
MoxyHd+Hodd9+mYE2xUYEEt6gwaboBGV7W1o+Nchfrsszwzto2Z4+VmE8hVUpQkNTt/lwrjYHaGJ
cOok2MNJqACFMHNOEDYAzZuGgFeEo+KOrkilyjwEHK6e2iqrniQ9/X8fnd7LLJRrdaxCMR43RqWm
VxoS+OWzg6izVibhivVZiAPl+aAVnDoASqOVH2TbmB4Y8ncV3YmlTtlQ3Xa/xlNXDrBUSTSkeVXX
PTo13pStJyBnWb5xBI5S7jD7g4vgd3+jU5YBXYBHs7CA2GW+m3MuQ6dfohOmnt2S10j3LAUQ7/iU
rJzAASmKLKhtHNDD5JRO+oJDn6Wtb9OaYkKEBxmPrEL7aX/3Uc34nW5dhBJ3U4x3hcwqta2xcJhb
YrJjTXaaX0c0GKMyadJHLBKvZUd7CR1q0u4fpLLn6lrYowU+M7u62oV5A/AX05E1482VJ+GrQ/gt
NSny84QuSN7rz/Werp+RPmELC0oi6mMz0pLbC51Yom0fHb6DuoyhczkZTTL8nMaEMfV/Ry+Zd9fJ
HgzWM3A1FS8+6kfPZFOTPIAE0/Yv+8Ifr0dS/uGK+rI2+OsGmVmGgeGiTGHxgaMVal4SBdJqH0ls
Oj3Lh4CWQdmXVDEqRC3s/bEZFKr5U8O6hLZnJgcaUExvX5g0VL/qEyc4VzQp04n0cqxQe9os8P5n
6YNG5qAPaL4qrhEDS3eQY8UCnzl7TP7ahF9sfcYYhxs7cBBzP4rwqole9gZWrcPvQKEVtRVB/6Fw
+CDjrU4ugbmaPj7Dwpfg4RgbrTFH+njiECpIBVcWlxOrSeCPRzKz0gcOyNIjb2qI2mjav/zZktKV
rwtaPOKhqabHjII7Uo0Q8xl5coQsq7WdfPaoGXNnA5qKoL1hDRtg85LVEtwZXMP7qE3uBtRF0shO
HKmVCEZbJC16mVq1OMiTfQ/zAvn2U6yns+MXfR1R4gExv81BuBA12h0q+slOQDG2FyWDmVYjJ0kL
2L99dY9iDkyHMY2wa8CpOubonzTX4WiHPCPOGtDQ8ynMWTBhgjLUHTsWr88ok/4WFQF70Z6DPqgB
MedHd8WD0Vl+z4oaTm/CTx6qZhzNZHN8SrDKpXDiuwaFw0WsUIDkSBC+qviO2cX4hiT8hZsTSUhY
k5erOFfn837/FRvfMiHxaruqQOBrf93C0njPi+PP0ATnN0DHGOZ8H3QblJhansbx43kP9OxS3NQ8
VIp6tSR2Kpx/hLAzMD361HpX8DiuBLwlmvI9aH9DZ1GLTbBB4VC2dpTAZYBa4GYBLzswhDhgj/sH
nokCk7Z87qms9KQsQzaNLF/Ud3MQ1iGdMpurxnSuPFOkoIpjmu6OIy89vBmEKcynI0iMLI8BxgIy
4U9cJMqJ0VfS/uHG3eu4EchSRvZIkEkclEM/SA78J2tgTxVbDRvYqCXw8MeL5NlCPgkClc4MT9Dn
4MUMvriPfwYDh3QsHguIItrBTCoHaA4yMMJbSaQr1tIMEJE35n0p3+qcs2Ez4ozL7RMgJenXQO5Q
Lz28oIsfTT/7FxOSqC74If4c31x18OwfyrDS9/VY6SoSl5l9yp4SneDtOar5Svhw7vUeUnGEwcew
9wJHZAha2P9Gico0KJ/XZJviYXjBVBZAi1/waTFfTqiyCoNTGso1ibVxtEAIIINDqEWh7Ctf58TA
b3fHU6GihgCzCY8YBZM9F9fq/Rca+wzTZHXUeLFA0bR8o/7jOXLZy7uWdHAwApLdaiIQE9b/33Zs
6ySDG0sRwOvWWsmTNasc9o4T9ASVHg70eHao5oF2Z8Yvd3/jdweFbXtjvUQFNWD0c5IDzovhnsQY
PZhsIcuIzGX9U2+GFiBX6R5W816iDeXxOnKgj2x/i5etaydhY502bDEaBYijcHEAMX9t/YU6FybM
xIH34LwGP1lU40hgX0e5cZ96y74zXTq0G0EiL5us4ajlcclfsv8cZn9D6zdIxzAI3gT4FT9sgOKK
Qu2+HEmBwmTzn1yTk2v6Lar5La97auLeWEVvi1mD7U7v7fKio5rGxnO7LDerOKjg3EvV8a9laV6G
6eqhgDthuSHg/SVeClR+vqzAJmj7rQv5fxPiRCqUu+san6BN/ZcSCNJZgBKLH3O63vAb70jSurcS
xqSdyjD6b+dJWX0td4A8ZeUaSv6IJbJuZSQAiZSa19veRowLWH7ub2ww7Vr+c6zEwm+/1nylsG5k
RVbr+Eri6xBO6V6X7RbZPyql3v/Ra/dXacgc26choA97g8EQsRM42M3627yF6ONqxB1/5WaMPcEk
U6ieBFrbLI4Nyh2Z8kRijxSItqFDGLWOsS7MCyjFtPEBjkZ0rT3VSkjRbtW1+XCeZRHE41qdIMfS
aXuj99E8EcORJnFxz42/cx6jLdwMLQCFCmZlFPKeOSYl56bYaIFEoOqejRqtkbrfXOajl1Hon/by
DbGbAXd308PgphDC3vfdZPmqgl4MgASJCwBijNV9IlUGDvgvQ+PtEZHll8J5l2DKkcNmdc6TOVE+
zJNNnDhfc5vNYvccIhMmsvpzQPQwGGKSK5ZakaM+Kg/HW2kFfip4VevWa5WGjdo3dMsevKrQ+xpP
zuA8aKE7uBFOmBQn76UdXh/5wJpkYHx4Sf0N6g2TpUtjbpSR385jisK6k7z7H9Il2k9cQ6a8RDAy
A3rfhvrn8oliAajhtQvmQpfOee9qR9O59h53HI2VKYteGkrnnPIanzybuww+xG/t6fAGv3fQXfHT
MF5Du1bVKQ52rlh6dZajRbL7lBLXkhZyoD2AvAg1qIJUAjf7+mx2z/sD9w9Hik21v0te5qkhK7sd
C3OaN20sLSlXRkYvmFCibHgH7dpCBb7e/YCvQ4gIGUDq8hlxHu/1SBb2UbFRaca03vQVvWgSCuYl
LmRzgD663/9IeN5+42t/xRPDtP7PkDihxEWy35qwEq6HlSA8QKIEfUASOYyU08Meqhhe3+yqFjjq
idAHub0hqwBDiz4Ki3f3VRCQXAuPWmRTkN3Y83LdRA8lO/QhbMTz/E2BHEkcFrXKgDqdNw0yk/wx
FKHdNcxSXSECYE3kOHzRxSUjr58nmDTsKGQjDH4IRI9Q+Cj+gSbgRCQpEAnPsrJUd35bW9sluDRq
fnVPNz8i9dTSZT3WL4N2dsIGb4vbsF/79G2tPBPb/0fQKssR/rM221PULsurfP/m7BPydbI0s0XG
aCoMZBmVzzTRXiwtthUoaDlLz+g4wwWK40G0I32NetcEbpAuo/YJkEffVHkXBBOB/lYo0OI0R3Xc
u7UCz46Ty4xvfgYFWSGvHDRcMLRc8Zx+LdHDsu+HojnpAdm5xNNu/j5TtffcP2Abrw8p7kflsPB8
u1PtzNgoofiN/4d7F6b+w4iN8JvnUEuqKN6QLRf/DmWp6UJXO3K71ojYxJim+E9+mmUykjTIpAZA
mkg1dR95uuVQ9TOR/n3Ga/T7tVAV/dRfiIqO7CfVr2NruWn5G+fiEBzDWwYBgz49nTaOC1+jOT8P
00oTej6J6Dr2sU2QOnM/bbwKMTit4FVZQSD+piTu/VAxoSs6wixHMgcLnGFsqTGkA4gQrQw/nNpi
Y+n26R47wRH0eZBQ+m8akTZDSo3gndDSx0FrBRMLup3flun23gqUFgu6noOMwJMKK7tV29AEe19b
LS8y+sQhrLPBvJs9jpIW+0/NPZ8ocyAODIQOVs7x7E+i40o/obneN3P2/2zu8RGh3joGfMeY99Oe
fqRXzGzkqegeFZwJMi2LQcVCthfKGbXP7GtWl5wtjww4cQwKYjaD+DtSOkgwkp9JLMKsNXgqvUhp
DRu00MsDH1AaYZzOmzHOt7gI9RVlT93FfvLuXhc0cubHNpW5YBwLGzzjcY2tGPFt4jMUcGUSQRIL
SvNfFUsAl4RF5sWjqltsuUBtJrPxz32BY+iJBzrxY4lteY2nC7FejeXlR4Wmdl/QZ4gPS0ImKUEV
mK4nMYWQU3nZVXzTwCHUx569weiAulqGL92pCxH0QTBtqxssbGlyHmFoUc+l8H+sFRGCITVvCYh5
wPXbF2l64jReO+PNQtVCYCtZQH94NbbRXHMgLZoUFUt0HjqHF7N7EiFf20WFzLteREYvio7UQuRr
RV7FLrgVDv8bsg5cMtUftLpcxXKvkqa4F1TFS+V0M+N6mNRAExvyNPgEzh7elKP452Hvv5XLLYJu
dlGNWUQoVX/h/S36pfdyNQDoJZEHTUtalFZtQmKcEV4qubmxTRKX68p/jD29x4HAiIajdFcxFn2g
bpA++l8BTgSFvAkbc2i5GmG8s1KY4QFIznuU/fn5U8Qq6bSiKTKENTj2qy1fOxXYXpv8msvNAkcX
2xCEvyxAjXkGkBKwxAsjTJ0G2buY7vBU8okTprjRc4uKfvV7HGTxcxKE3M0JB+WDpni4z5B9dPQ7
JwOAFKc9Wo+UtD6twxzt/WQgxUdBZE6yqsgAnOLesFjrPbIHaThiu85Pbq7KmbtWoR84s7g3k0Tt
2IbY4HbFv/uIdKYscEILMz3aQulzXK9VpfmQmWZdN/c2Y5xdwuEQI5NY81kV51zAIyOuz5X132Yj
haULWDFzVgI9Q3preI+6NQ3oLrBps3cf1yt0ZuS+lZUekTAdm0fnhfWIXzUArtLvV5K1g4H3yucg
SroXkHUPej/CcsAms3v2Pxn0nThVarbBloT+QrEVkhx8GizH24L2ia69N/shhDwsdQwIoB6MK5ea
r4REPDaq4bW+SWh30QsVAycRUN6wBbbbEmE7w79+wAWgCP6CCwSn5WBAkTEj6JgPJxAD/yoKRFzw
+fSyeCZeufs1Q0rH6TFqJuJ/8aZoE0SorD5x6aOOc6GQ0LW2CDPz0+nx5s9yG3wOvdGlZaivBXjw
K3FGEewLy+mentsioAjD7GrPvA9OXb/pAVao9oqHSA6OwkmTrjOJHt0VioQTTreXfvfpiApYRzTq
G8YoX79H44VFKJSXowVgmEC8RJizYHmxV40Kh+FGuVz2c7EmL+YajQWQYVY//ntQPSOys/jHaLH5
ZdYbdxMm1u/QoLDmI5Ow77YTiJoeUktEyf/EihZC7XxTWK7JuaqvPov6vZ2d6OYDZX3YKkXNMPtF
flWM3wnS+WkEfx0ZyATMoHu5Cj2nAgaFynXF9WoWm4ZXbwXG9bDNxMuGCJneDavM+guZ1xJd2OFD
ZeS5kOxQPOnEIoCKoYmhsVllW8eHP3+694dZNFD1vaLoxD+oPNYHu9zr0065BBHA++JZDRT9M3r8
Y1bg189TpVggNTX0w1d4wjppd/pHLMMfljf9CeHo/Iv+8esYmhVajYdjCkeouJBQinzODF7ElXO3
hrwIZrgYm7hkFAyj38P/9lbYycA0dAJMgYQJ1vBdvIJPBCE0YCxMsZHF3kcbGHKKLJ7DZig1sRy+
lHjvIUPUEk0/fyc=
`pragma protect end_protected
