`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J+LLxG0D5JxlyKEJjlDLJW0zyT2TumGrunJ/UWQaAdPyxunIFDyryQ/iDZkYmQ4N
L9nYHIkAHi8vLFhen0efO1UBsZwXHu4tvf5HThmvU5oXSPvKHFuJqP0ZxjhvUuvx
qfLGw3O/Cj5Ait4ktyOglFZmmR3fCRb9Gkm35NNLPi4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6352)
WCu7U4rhehvu4qnXMYKbxOc11GGXOgcjs+9EmoV5HJbm3z12e5HpgvyMYqLYGVve
PS0o5iFRh+k1nHI1w69PkbdQu270PRHAw6XsdgBvvbjcPjJVQp4QPg3f2dClkwTc
0YfCBkaW5p/LbUEkltLsDcrJm0g1TRY6jbLw18CsiHF5ZF+4YjcwMu6WZo9/rme0
GJ1zERRsZ2SYrvOyGnP3PUNjbCj5HMMufQzMR2lX61ayEUXJPci8CO9MI913WE7h
TNqgdw1CX62qHACrGzLEP0qrGPvsLKfluFOTUjxv5u26+dtrSrBHgp8mzhrMd7af
mo4FeRTiUKi3JaCucRe6aY8hSY74Rpdwyh2Z96JCQOjGVvMJGOD0Kw647Qus9h4G
hynAwv7TsXAp4lwFg+fUPaH5soX0Xlz/qCDg0gkla6YkM91eNNiY6jofJZAMwz7m
fl9iWW1H/bNTLICT3FXYJ87Dl17v0R+/dc9imqjuU24nHJZD6MXRufaFPMi5gsIX
3OWNC0K7l7N5FFNdfGZjo7EBXHilYh5cGuZrBAAl58Zwty1Zp/RaT7jbhxEslfTr
y/nHGIVSi99bePdA6Qg40tPdqhrcpykrdsyBnUBnchyc/TrWyK5NUoctXMSnfPTQ
OT3yiIBzwDHRADE7XzbdwWj8vBC4EtkOQI54uGgF/3BgRac8VdIRsmm1KfldMEhX
yym9ox3BLUIun7ErmJHJrtikgM03SZUPbnElIq3PdS25WlLr4cCwAkXS+OwczYxo
qe+nbHuqWSlAoUaLkmWAvY+GFFBjxmMe761qYWQCfHg5zwt/3/ot/XFrZI1H/Ip7
s0FsF5vOEqakY07unk+wrn4nYJqAJ3jmg6e52GBkgwZKjI6Maz5tfMIZHnUp967f
StcVfDtcHw0JVCFd8dwPqxQwuxDhJdS93YJwiHTlowI+HMGquHZ/96XIM1ziiRiS
xHw94RZpUF0clLVgeFBdZhf7gIxSLHMr/mzCG0f0KajkldGHuBiLj3AjGJKDbstt
H/d/ZGKcupHwiXvfd4Qsvgio94kvXcABB2u/WUtGQXmCrRhJ7uqvvhLJlj4TFsHE
zLlp7BHdF6YuMvhE2NqgtX/XZMrxB1m9ADkDvxbYaSA9Baqs34zCBk9g+NwZIOxJ
C4ynubqS9bp6GCU/ES4lli98nZywCVRivDhDsIZkDJfdAikFZbwaXQLGD/z/jH1W
IKYT8zivuPx0rmf3OPwIfEwIgVKxOGmhi+XSjTpC+Feyb1zyf6O52dyFpF81mE37
Fv6r8wjfJxu1jWgSzHNcZZ8DdOrreVRsLaUD+qTfD0kN2ZE/cVpP582mwJBsiBDO
mT95IDP9vqsme960UcZzms7Fb5B6nqN+Gi9RzD5sEye4lcLJCFnJaJ/fTiEYT1UY
YqgIGw+zELa/ix7IsWEBjsxNlST2dCuvtxtIvQVM11sLKj/aZAl6zojfENFendVD
wY/KGJ4qofgDhqQkYys5GIH9DuNCVrFa467r33G1iutyeRqS/njPz7Kh6aUNdPLB
bi05Ic+Ghba18lcrTZZWM00WImVVB3qBQGxUEfQ/1Bf/r0iWFB/k4A+cqGRFnwM2
E38Q80BFvSeKc0snBbUuJK9iMw/fA2qZKqXZsuSehJ2H4d7sUNx4AVbsd2X9/8lu
OUkbFqFWO+ZEcUOvdFHojsPtCub37iQrUUrZZkTVAvsWtQQmbOc7r41C8g9uDwKH
LCXiT/9UVeC7eeYrflhOEfQiNrcDwlFXFgBROAJxZnEc/GDzs5TGwn3GJ+t1siw+
UWJhyJtGcVyhoGo/9oNWRQ+e91YUmwXfeZENBC1je0N7fW48o3utv4jV+CAng9iG
YPiu4Xu3twEVmStVbI60MpRRVfObTxmz5p7kYNG3xaZjH5LIqdc/IUnr/S37rvov
wKM6M9QeeN09az8HkjryXu1hyNefMEM+axCbS5QQnuc3xFJpF+g+GNVIS4oSE0bN
EugtSeZkRyRCbaSRBj5OReR+62GcNy0kNS+G4vPjm6MMc17CM0aNRJZEL9nM9Zzm
ETpujp9mVL456Lmij6nCRiNSD/Ouqd+v4YrsnpDmsDBSHe0cTwWdSRvuNuU7KUDs
fL23oe4Lp9GJboJI5X2eVUW+2imLhfM0MLwYz/c6HCh9yMNtesqivC0DVlENma5m
8IU9ZYqkN1T02wCH1oEBmPpxYhBRrBUtbGe1syofXBXsWAKRGZ5vaKRQQXe4tUoh
IOSju1YnvBdZMLlCXSga6FmneCshXCRnlZ7RISP9+5sETeoq64wa2t8nu3Bn6kgO
6lG1N3msGrAGuuM9w++DW7yG+Ts99z08P2x3+j9t5cZPIDAbrPVsuBc/jm78BBVb
PtGoopVzcAwwQjVYHPuUe1xHFqHDhDmkJ79MOwltSezLO+g55GgGOlS4fhAczqEu
SdqcAtaNADuyX7Kced0hL2qNq7Xjz99LS7mbx8l5ROcwMuE8ZZsdnozxMEVrQC6P
11uuSK3e9cWsahizO1+jdpoaFxraKuJzP384a+f9MMuv/NFIZ+YN+qCAwUZjO9Ra
5fJMerslcM0QxUNSLB1X64RZFvjDawcWakcDxCZzEPhq32elb+sd1C+wSLjx02DQ
03kGXorkBRNSX2CzzuzDqARE4gn75SybxH5ragKxi9iebP1Ryj2La83RgO66uwyU
yNRM+1f8xl48h9FeRTRG/hyY61XtW39p+vBkkGau+bxKS9RJyJeP2ZwyLCcntyeJ
M3qBmOcSywYyqG/2N/W0Zcgsgm5kCXrfESYNAgz73WHjohufyq3bxT9hlxqXvk8O
8jFwjVGRJAqOzP+OCE5MWxi6AuMsHmzap6QBJIHrlPBJQ2RclIT1wJs0rKHGQXoN
WbugGgRuDrAMcW8nbUIfnCnaMNa1fAUBzjlU/Xtkzrf9i1eF3GLd187kDwT+gYVd
fRWpkNz9/8aknQIEzkOomj6o0JD+y7LgA9ispvfymqIr2nVzMsuHOUw2bef7TQGO
JldX5L4iniGvFqAoKQTqV5sykEqii7B7qqS8YaiIM1alWC8TS3O8omeIQzN7MQ2L
9MVBo4TA3/ATI4PSsRYg5smarEzLhqpUHQac6JQiTIlbHLLwRjPk49Q8LgG5kBFn
97zxkN2poVZ4B13FxmJLU7f8g6DFo9hPLcD8nbbqRXnDXEza0If952yNgdyW4QPn
HKxrvBn2LjithhmP/yAcDWTnfzMk10KBFSMMRnulcF5jg8KuQMNiSsmpRWHXY+Nt
gITN0A1JSzu5LeJ91UBEvZWZIeZ7UAEYLivOoITWXTKclu1JJCP1ofW+2+djQ1pN
3CjO6vHXHEdinkOBcPKvCYUBWl8hHO7PokFQfZ7zRG6z4eS3RKbHaSeF4xvcLD1P
FJ2PKc4484zVdAnHpCj8Ss7QI3zAHyLdeiO8n8Ujpa94prPetuRk2yAXBBBf2wrV
p56Kyi1xQuiQn5j9XzUQ8LhV2iBxEekEIbj7N0m8GQQInQfjRckUbTyKlwfADBZz
5lsdkIO/U1NDV6MjWSCoDoqJ8MyDpLvkHD/5syWPGbyUBiiD22Ixj7IAzDGxGCw0
ijHcw5ph3Si0AChFB219wlExchymPmXXG4Ploo98SFfsNS8cLkr7cdcyWzIs4bwG
6sdHshL7f0eF465hOBIgPiWeU6gq2YUHf8XFm7jtHOnN7N6HoG7UnDWW+d9r+k7q
n0N4RlQId/id/qoos2l+hf9JQBj10Ws+2ZDjGla4UBN+8Ov5/aW0KqDZGZkZa/b1
AWp8I6IvY5UuQdXkRemIZPMcAL+t7FmgIs3KxYcXt5mKR968Ibs83LpnEYhSs6s6
agm9Pif+6iBHnnpQELxLDdmCPeG5jINpidmfZgPJ531dj8334+rlKHWsOKVgYCpS
ujpX8fw5xkcfEUbba9pGM/voyoW+6q5jjyBqAa5c/08Z52gJHRtj8kUbm8AE2ebi
Puq3qvsmtz+35fU+FHApEU3B6ZngR2oyHgBlZe4w6uiCePJ839fR72bJBWAkT3GQ
YDlREFv4Wd4vhBQf909RJ7pBNjFov6gaKBT9bah9FObU5Y/nHGkCJinxIp/pmsFO
JYik+XP5SE2qKjNEw/gBRd2K+Py3vzQSBAexIdk/1gHGtk5h3gD4eIeAlA1FSQwn
jwMnvRLrJHoSaNitb3o2aWgyfXUTuSK6Y0/5rUkE6x6ITqQwRegwma+QKtNN0amN
BuDfhPWVlI4rz3YjqW9ocJ+Xr8rKi8Q+KSlsnh59Mpe6I0kmwTYAtEhRSCE0J8TB
M07IdJHdTpOsUpC3wtqXAqcmUOsdpO4fuDd6UarzwVRVEltvhJl+wJp66oJ6FQUy
O8yaxM8hYkQ5Qw+VEPqRHVCntcQp/DAB03lpsTwXg84CzXlcpjasA/PZE5tUWBNz
LB0NVmy7ymarFWKNvQGSJfAfV9No7AFQkEhOuujbZJqecNZudFmUEMZL9qsvNC8P
1qKTH4Y01hjgGO28JZN96gO2aUWYQRk91f+B6Hh4FkTS8kxt3cuRlNNrwLFxvIdS
mRUpqEGRfsc8xHcMTWah/+TeLlBd9XQxh38QvDdfNUq1vcezfDXlcNriOBj4zNCr
lEqKLcnDnyFVCD4OFELA+5nsUSWYjOoGCMPMlKgANXWTxjNE4Ccxivxroc6qy3sG
UPYZ5LjyGUXI1fKowpGqz/7WTjP1R3ohjhRsSRMVQEVFdIDN3EZZWOvRXDr/BgP1
aidr315kTRlfC5ZsTlz4ncaN6kAls7nWLl2DzLezAfZSgDLtuwCur6bZl+JaFwMk
r18KDfT/VlDl/emwohlfXzD4WxeA4xDVxkOAJgkZKEHK1ujR9AaKqTRB9DW8QEgy
62uvvEZtyOI9XEhjnuB1fCxlkD0TklTWsuJ7ZGcy5MDc6T6rvTHFv6y6ErhhZsoi
6yXekiHDRjVWO9Fjo4068OestqcA3tRdqs6gsAiAxqA1FwdNoxDuyLc8XxTcpseQ
D5EwaZFRcSeB4wj+xEHGUi1YcSXiUlZZZrThbjk38P43VqUCLwjAqmp6T6DaHjYm
e8O8Kj0Ty87mB2I6+gYbcdXzUAWafSi0Re0FZ/6btI7adc4AODWlO3wfrsJqjIqH
6zHs/rkiLJ3tUqmAc9CbmPc0UN4ZDwMPcS7IcFZKmOLOjOWEo2SibcxKdXdtxG7c
7ujpwRIIH3DbHMwjSNn4d/W/uNR1nqMy4ez6l2g+kXL9YallxULOCp+8jo0gKj5T
tmxcw2NCt5FhgHs7yqtINa6R3OOTzTjOZaP5kdvY+P/5kcai9GJiKAYVQhEMQDTE
B4t/5JwJQiNwRhkP5MHC3kCwlyTZFvB/w9/ba6hxdLA2o0/3yCJ+fPvTUdfRpHN/
3NuGxxH+ssSVJJ7YqbqKrXuXX6aA1ZfN5HaHeopzHqWIZhtU+5uxA5yl34hzcLPO
bAjJ6tQtAEURC4TFv3hfMHnRSICiOeHmfzadSzPNsj1IjQ/l8i+d7MzRov/XBJun
e+5R7Gcn/FMmOhceDA/fVKIOdzCKHeueuB07QiNVWmsbxqImXG/h1cZSvessPCju
luZR5IqDhyhnslF0emYodjw3812+DgJ0USmNw5a3nn/6l4TYR+2GpsEymPcMtJ/x
SrpMZIJPmDBDVf9Zlz5P26DYW3eWGHBM0E4FCCN7ar/kCpuBUZgj4zk/HDbQBuOJ
FOO66fNjgyY2XLieiI87F7OuuLqMthJNRyDzSsYhrpq0D04WUof9wyAH0U43a7I+
/wYnZXdOPpbFDOyqJl/ljzhe1C9mlfdLnhNKOmJ8ZjWnYa5j4x8rQH+C4x5alDlO
uQhE8yMjzRAodvByCGq7HpHJWyHghEwQV60L042vfNxgZfq2XDNYCBUUtQF9Xe7E
NvJ6Su4rXElmK/mT2jsNEa2mbi0B8e92t8xYEsYqoxOWToNWPfd4AILKOWRxGxvt
QX8kNFeWSaQkg8cqgEbOx6y7Mq/hioKh7oa8l22GHyOoyFVsQ1kexISKBI/PAwAD
sz+/1yzFdQNnS50bXCliuGC7KKBrjGo2emUkSfzjS4hnbli0TikMcuyYm0T8Ozs7
1gM5nrr5TCuRT6Mygz64Oeiv7wOKsX3ctRG79a+3Bp+VUsClfNPmfJEh3kV7lWS5
CMGLTdhZfYJMxFnrupzG1+hqj+rCgH+eh+lteALvU5gv9G2w4UiL4Pgfc5f6gX7s
FCOz9YgYP4yfK3Rdu7+ZCvbG6S/8ugQygSPIGyTezzOXwlUyhbBl1GrpHa4emfa+
PURAuaxysitQZW1dyDRjbkWWA2D5S5O3HNlNoVj5qym5ylmHpurHUix56H4F8HLE
BURtjmfR7fbkdv2D0pga6c3sekK6HNOOogHWLEW5EN7ixWGyANCMhMorFvw48U3u
OX0wl5oMN9oGBz1D4imM8b2a8BDCuYfln3il42aiSkzVRPKd/mZuNBr97KThRB8A
KIvzUOX17zZGFXRFKFO/l5tG394dESYWqG6PpWR7FbXzAC/HUZ2Ce/T4tb92BVhj
QZd0cqlbIehRrfqZics9NRl0EqiFKl/qGNhMmDtvKgQXrlKsJlYRqgEaW7slZobJ
MG6fc6GZt0k8Yxp8tL9nzU/0tMb+wiV37/cR0/izYmgV8mr0WzaP/sXeFq4uI1+4
X9NEx6oWtPbZWqvKs7jBgh3rva+sHx0tfXiGgI7tB+U+0r8y/N/hyhJUYQDiHNrR
eC14hOjLxcZGBDKwwrMEtTEXukeMjGjbXRgu3ptLFHogQ7XK2e1yySLcFoNbewZb
eNrVgS0Ta2V1cjv7795gZvrk9OAsEr1siewKwqnDBKyZaGmC0I75sJFPWyizQgFm
3nivBu5kmEW2hyAmzMDA7lFNugM+0rU6KGc1eFvYjwWiJe7g5xqZiQc8Lt9JhvAl
KY6Y8mvAYJO4vunpAb+x4xo7Luf4dKUbnY9CTvEHHxV+T7Ppw6zALfE6EmOYye58
SOO1nnvIQj3/RL7DaEL3u4f1bNgb5TDXVDn54rNge5ghcgL85g9gq83akD0h3W95
m8GefIM5VQPD+asNBnUVUHBIfjLA5ebv8EcazZ37u0gvALCy9qvi1Edgm9GmeAMX
JMcTURUX308YwHhtiflGvqQVMuXhk4bXiHKxqp3XIb0LEUIoCuVFmNkcU82chUHj
LnlwD9raifMZyrZISmm92zmuzeAukOhhiyoGqn2xhBMWeP7yNrSsqBArB7lqjZTD
d5HAECj8B2ly5udQzTotKigsQarQ6bWFmQIab49FpGkigQHe0IYPqsfjnmbPQkDV
KMwOlZ4y/lqhdpjxmbKL/dmG/AJ2/wdExgKgdVqKMmWDy/vgphqpzreo1KjgQv5c
/Om5Ik6sCUDzEXT4tSYxswWNIEpxWxYucFJ7S+UrAF/pxmD5fLe01IH2Zn5z/IPI
24l+/abOTLcBiJ89VABmPG5gdAzzoH8cijcMv2MTTvtmdRX8SivVz/tnBuC8FrOO
7C0nNr3SRvZ74GL2nrf2ZqK1oOZ7+2k8+Ny7TcYs4WOpRsyK69UVGFg5OWP5mvnb
AlY6x79AZWHdnYgofV8FBhpIXzONRcAMUyCiR4kJ+BwIMCI/UyAMSScCgWvUO5UW
bDKuuaDaofRjLKnxa8f/2i1mgYhskhzDLhoY1LMoKJQ87hFX+JI+XQcSkgmz+WTJ
WFkqlj5mcm0EB42w1A185M2eAf0WsV+9TfS3jlXm2t6FtPuKd42trT5HdTjaGuId
exJq0FRB8OGITPMOUUQQaAPRFl40kRfxyPX1gbmnq37uev6CJ1kkU+kwFnzaAfax
GU6mhwe6OSHSO6PM3sApnAQUGA+nuyfn4Yl9+ANSaFgfatb5nHLquI30jqYf6H6s
Ek/4udwI1LZdVtd2HJH3rvJssWIciSlc6zMYvefRDNUJYs+js7bGaLSWCCDZwHU/
dYUvQqM9uKGyDNQ/eZctXRrZXclUkZA+ekkoKHuK60KIqwCw4oM0m1QUZe8SGKjw
DqsDmJCJTqp3h+2kTMGzdbO+G/ery7dO8gsby4tVqiJufLjY3APeQa9rTnghr9qC
5EFgLB7EeW0UAxjlnDKd/f6cV9s408N9sE+tn/8qOtRTTBsKBWhFbdfPuMPiAFwz
5ByVN7ltD1/Ct68nwaaQpllAiiuqBzrcS4/fl3hw6PI6JRW+a4KK63DxzJDwWMhx
yQawwultfOjaKRG23EUdvBpXBC7SyUXxtxpE3ma2X2ZH9bKwUL8ZgJAmOWEXx7E7
mbYv1/cGd5YtZs+T3PMdYMGRaiwU0Ccl6rOnVv52N8skPWNwiMuUChA3xlCuVXf0
Nk3/A9vCd7ELCN1kqC57d6f9Wa+GSBpSeE+hsyIkMhDv20LavSm7xqhROVpHQ+9E
GyV1uaK2EaMe81nq1GPu+DpxIZEHWYSTWWyB0fbnIhtjJmHSXWxXsrwLDyq3Cr50
mdX9PQ886akFvSIiNhGoig==
`pragma protect end_protected
