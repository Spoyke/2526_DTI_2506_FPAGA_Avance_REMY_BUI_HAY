// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
p6vhehpSCzmky2cBqwiUIvn8Tu3W74hsqwFy53BJcnJUY7y+RJlt9AILFkajYZrJSChOB4m6+MBO
LPh/h6YXcAYS6UyR6nCZ+qNA38EznLK6uAO9OcaRbEomUaOegqk4cYRqbo3YNFB7ZpzVYBAA1KRi
dKhCVPft8gx0F2pXp/PYbISxb0rnVg7ZNU4tRGxOPfeKSm2WPRvoqohYkiF7YHPsC/0qOjjzHptp
DHT1WYa3N+C/+/8VBMqP+j+evwpuxg4OI1OrZijgmJaLiMjLP3p8M/7XAUJWB8DAnwOWhxDY5BAU
w3VNbo0nKv0vomNS1135oy8+Hve0990cVNPFvQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6272)
qcoS4VUDYzmj6W+ypA+wjmlj7Xrx5ZJq6w/vCGR+2L9V3m6UnEEeh257YL/5IXEij+OuiunHVfBs
lPE0Hkzee2Cmv99Qg8wf+r071Ml7NcXs+Sq5iNB/5DCX1300torFO388LuCLptE757bIVZc+GsUG
d4I4s+gQgq0nAez1ZWew0pFEr4q520OpXBxsI2EYdx1q0a2pwHT8/PqnX0tG8FWHlWGMn5i64moV
gSfE8ukjdWrlKJ8qY0a4Hcrd6ABl6rlHCqsgi82H+eYIsnxCO9ehd/Au8thPuZgb9s/wOzUkW/vg
0WhJbJaXtINsMI/NvhRtHmJ2pYk19cJn2jfNrKLL2M1ZOLnjBbbOj2U+yk3KIR6ooqd25F1rVCWo
hagCREpHueuIs6fGCRFYuf11KLjiJIsKWBoqT5F/nQQtsXmg/L9HnPpIv9PjfhH0cB5cqsDkYlA0
bMoIzVWUZv71PWHPMUPLtPYwZqWAjZrjY/REBxobiQtez5JJKdMxLy0JGI0ypTANwwajXjeUmWXD
XGl2Ge5zTi5+pSxTKY4kuHNN+HcOQ76EUC4CwqdSYbPYBLqGDuoil2/gEbpIi97eW8AnfWTCrdqL
qvA8xNGqofaqgUGMgXK9D9SrNktk8AjD6FghL0mg6cmq5a+chv421zve4mIECXaXlm1B+F65Oyfp
SUl0OK2jNRb7tlctVQ1YQW83QZ2tX71k8KyWpw4TXZVX8YahljoExHTy67tR0E8tT4MQi4nc6Ckn
pClQ20KMpTl4EjptQfrlpy23Sw882Mp1z4kTjkR3hyl7Sxq3qj2Hi84Jxo8w4ljKg5D+lFNDW5YV
e5wJ4V1UQm6Jp2WGOWVHwMo9hiBwWoI6t4xNA+3i2gBgYZFJU6sz6UdlCa4/eDPcVB0nVSf0WKB/
/bhi8Q61lzO+vuCRzCWHexiYh/OxSlqxtxu57kjTzSWtYtT4tkj2srMYNcQJsb8WfwPwjCEZNS5R
5pks+pT7GvYqbCMyTky5mMbDvPGgAoD/49y7NrOU/GZPGJzIEj6UVsIO6J1mUll6NwguYXRQ+wcX
mPiM8+SA9D+qjYNxOUNP1YAyum1sQ5uttwWWuGDg9gYBmbt9Xv5nGX/TMUW82l4tOLghBchw/7MK
7BcBe5T4nsXaPWJqcX/Cj/M3ekRUSEmJchrkQV1Ynu98pEE8n+x365Qlt7j/TPS730F+f/WVgjTq
krZF1nTElAuqjv8BlP/xqD/rUKzzqgyhxMhaS+5V7ZJeKafpz2JW33y9lj7iORfxCHDmFk+D3zo8
0qdMVbpwnETg/0cMaraT2IucmMrSvjV6CMDNkTcC29k3euqpLliEhcru1o+xwsDK4TmeYue5PMfz
YVUpv02qDvkpJSmt9QvQSClQ9sYwZYMNkqUW7r3naAeYQKc8IjW8WPhENn3+mnnYtBNzJI8hwoig
Ce0Jnf1O1vk/1BSy1XTjYKZZjnJxLbVOm8iAKhEW0hJKCABBwTyXMm04sK8Yo2y/9/PHd6O6UQNa
xVcCv3ybj7bZHuFnJ1oatuNSAguo67NRB8Pu1T+tOBbLh52t5Dm6C6KSnfiIcYMcQPuQNzmRADi8
DY//0807cZFpuF1C1J8tB0f/U431TofoxTwCuO8iYiJ4P2nbdUs9OxaXjTZVSx0Fk83DVh74Ywt8
05q8HWBTthQLeH6/q/4nt9G34yzl3xL+RIjeSYJ2wf5/C2YIwCQxLOilHkPh6eLIgOUhmNs1mO6U
9jc4GbQ+i+775FrlSyz59/31eLG2Fog2xo7McbB0/CCkXU6ioykAki6Qk0GBX3wwMwpjhMsPSnD1
kyDxUrmWvrZYEDsRLwtRNygcyY2wZYGPnw1k0Uuft8+NVJaafrQUZK//G15lO+wH7F7iS9QUNs21
7cMa+sKqmfrFLAF1z0GYGe5d6Y+hyKmCcwmFeHyAc78FgnQLJBUvBxIUBy3Ha1lVZT07q7Rwtdqv
BsLGv7V0lCfLaXME2LdaE30/9dwVVw3iPs2QveApU5jfr+z4YZ3UtuZswNKIOJ8R/ob0WU4DRha+
TfnFwcbM8OmTBom9+ze5YGVDBSaPD4aiWTP1+mlAzOpE3QoMkZhrYz/otsu0UxzHfNv/es04mPsl
cATVcTl91IVy1pQQNttZBQUDtAKXG1V13GlB+km8Oyr9RRsOnizokLW/pRFC9UE6Oqrje4rjk1m+
MoqWTCbnynTe0BvXXAsGxQ2oIvbCLky2QMtWKbntKkrBLnD+hwplc2EDeyd4mfkTVcPjdazJ3+Rt
yT1QgHRR9mN42rJelyFqxJ79dq8vPxMIXFMstQ7o1iAxtuxB2neo8tDalYJjQq6zq9mvunftaUsH
VwDHtW8+PmoKg3LQEuVvYkkXQ+f6ELNJPoAdKSrHMSB4GnQcDf1veTZkDfI5+N13De7BIFxV6UY/
gUTy5txeHYlDwGgQDuq+isHhFgwTnoIV3aCNGBtGbAG9Gvt4aI+O9/Yjp3j3bE5EtGtSO2DHb/yW
PT5HhdbekELCj51TGUjWPC99rfbeOhRHhjBtBPSm/GLQUrzXDhJG6GWD4NaG9vn/724AY1/zn/D1
3RMjsrJz2q8UP/ae+IspziVHXPstKB8lTLLREzvkDNbhEejSkrXnyds+WK4Xrb8QqygHvYP1lKc+
7Xb9Mh4NDKE8GKbEBu1jwvpc5ZI6owITb+uQiiBDNfdmDklgKSLcQZ71CQkOT+KwOOSnC40254bA
Km9CmghPXqvICCZX6mDpFDBAF6EBcM2dFHqIsisAgXNokRzVMOnTCQNNUh7xQAetLwyXWSSC7DOq
YeEoTwIr9cDp8X3A4HOQgT3NrSPKoFSP8ZIB8vqNvPiXcVpVK2NqpwDLhzXWdFMTMEcXbj0t0hjN
zOLiiw/eRrzjGbuLj1aIk1frF/882t0c1rYbsD9PcB4XeJD8cLeWTzjSiPeROjmFUOkM6UbwEVWC
YIG5f/JBLnw/EoTKm2PnWhXkK4sFgAylZk4e9HUgYFORKAS7xMlcbBonvid1DQS0s3WDEwzMzPod
6eYHAKQEvfurjZKiWUIkdWoGAISyO57vXuXeYaETigYn5OOwmLNXVm+w+5ofLLfZLVGr0kKfQqkk
OvRBHuV0uKg9WRU/cYFAbFvuLsdmh0CQZkiQYM1AeqsMjOwno3b1ldheyYAwawVi6nH49tXj7cvm
UHG100onC6xc1UM7rsjY06xtcn9+mDQkIfo3VKLb/JzKederbWRHx73vDYX8djdE/4cCKLj0orOo
ClOiCCVtmri9jrU0/vzE+sy+pninXedaBoAVGfLW1u/JrPa2SEPiX/fc1S9xs5nmAZnEFNeqmt0W
KcrjLQijoUGphygYJeTqc+IAth0NIC+at2AADa9AHBnSYWNbuwiC7IFPuoEZY/qMgumU7RRzgLBx
mKyvCUUbVIN0MQEBS/I3loqdDo3/RE9oU1xgcPV3dGzZDODM8hFRjrtZunFNZ15AEwIBWLJUq/En
1eJPc5wzPWMjjiejzdFaV87MuowcGkwgGiKgz7F7/gz4pPuiJ/rmd3A3j2LfdZDmudu5FzxzzDkS
uQ5ZnjmgcinlyzsADHGhQa+/mDuT9v4GwhSKhdae+LZF4jOyJ+tma7TlVTNTopFb2hW7eeiLgsuH
3NotGAKaLOsJzsYRShYMgto80CGySVAeQhAApoFU6rY66TPLETrdmS/QhxWm/8wlkFdHmDxD0Jph
U9RtfzgBOxf4je3PfsKOhNh5pw5GYdeZO+3SvLG+Oa0O+iZ2IjuSSg7fya71ugAgQuFabbu9ghyG
qpjNSWbCGRl1oCr2iHhh3WS3GQ837EvlzhCSFyH9gLZJgOVuro7zzo+PSrOcntx2tY0hslm0ojh4
RfLUvXzUv6SHfWmCIwajDBqQYkK4FkF25Mnb1R01lB/UYBh4WDCAIUVfumHRJFxK9qvgh0bZfSP8
Zb7FAa8lLCx3Mett2wbSKV4vx7SZ11W38b9Qgj5RksfGzfmsMkLvQyxY+DBpqtDISmb800TW0EDd
BdUTOeYLmLjUKtUbck9KdoBHcy2HVlMBZ1IQ3YKBQddo0o6PO585K3h7h79XYwYSe1ZNvbbVbOY6
fLnxKOuNrMtgomeI3I3U1pFaPZXiTv6qFh06pAioKIXgvWCKwEZudK3JGPil1ICDCUQwnLvloHtE
egWu88s5p2FtIE0gmB4GB0KiAksF+Wf4KV5F5U3OQ7i2qc4FvCJs6e5JSWAzaGmJDFjo9RYSm47R
nrH+EQXJFaeMnDYfLbNgvJtcYUiUsOLjuSqzZBRjfhR3Iqp9bfd0QPGcs/RAA5S8PdiLVX5Uxf2Q
jJT1EMrgjkEluGrEtLAcD6edHthozsVKTH7EnFwz4TzdZlYNOgFw+G09kZ/sf39jGj2ohRJD6BWL
QwZl8/wVJS16le2QqLENGk7DqILIEON2FvcBCY65OzZbyvrFYxUP6woUYoKohd4wMspsIs4h0uzo
vyUW9cyCraSQDOTqEFkq/wYcMsBgC6aD/EC5VR8XWM6+Y0Mw5tsihXgEant2SJ4wKUlmq9kwub5b
FGbEiyxPF6hIAh2UXVLoXMja8EmiGxDj9LIurLIxpW7z0o7lpvpRhLsQGLYHKCj6LJ+fNus87kjq
xo8/r0GBK2sVHY5dP1ACPDMR0P46dnO8J+XLhxqmJT/p4PzqMQ29U/Hrm2KGcccwK2oGt+H9LNu1
8+FJleXCVs7jxKL46DmScZhqeKxWj4p8U4fZxE0GPfOUQiykkHSA4fbrIlB2KMBp4qmh/66zJu5z
0iTSmxHocN/9yGva7z5uMimQpyu3RPBYd60hsWiWDwc9nwFsNFwed1lNWKmYgFwYA1DPe8eq6iR9
AmZGBt6Ia7SifZVRorlMSfW26yarE8OYlA/YC7SOWp9jz66CyP6CJya5owQBNGiUpr4L4qqMUVVu
II4PkTcyGJ30c6H3/a1DYYnv9OMaEFiiNfvcuXJVbsA4BRnca0g7G5banSQGGdA05vlH1kDZbouC
CGbfJKu0KbKy+/4JIwQ/Zbkzk1eOLx8bIir+w5AflVMBpHis0P++tPgt+l8wnyuzvksg3Jy4+vgJ
pmxrA7JHb1BMk/hy4i1sauLRfC5Wc2oSdDpgxBW8XoHN1jAf/QJSPX5zjdlX/OH4FsYQCMHXKTJt
xxapfzJ/va07jTWrdkRSAeWR87WqkCdmO/gXE+gRp6+pAAKF/Of2EqOVxHRVXMH6lU/17XjK8HkT
UlHijhMAOVZF6KEe25xjq9pYlg3gre7jJauE7gx21jX0oP7BeEbMQrEkxSBQssqMkWDuLPvQq/j8
aZI6CNO5LYTfTpCxXXz7rl8YUuMIvAwhoScEejuqqFxIJCNRG793IHI9nKprxRS2kbyum97EHf7/
/pEriJMosaz1EooA4x+vZ2Aa1gQMsJl6+z25RdfF4wybgmMeiLZWaAhLj/Mncm8cMcUNoamhChJe
gaNuERN+IJCV3gqlKcPcU5HZMiCByK1yoRmhJWpj6e3jqLK9GtxwXh7L+orRxFxX6CskW9Z8tVHN
cjII3zZWU40RvH3Oux91lgJ0JcYEcS2hrUwVOrV3dSv42BiMrOXOg7ebKIgQ2nFAwb1cZ+izbqhK
hHZqLU/VsOwlb0PVhLB9s07N7UKaeOCTnw2qhJiI37t53HbposAuZmyQ2oUpJIqDaA+ehKqhOr23
/ceUQIhd8gOs+jy+5Rmvsd14AVUlhdQGXTQzqz+HICi1zNzeQGMY0vdwgTDBxeQE54seerfaIuni
fiuSIRpcMGGtWuxT90SgZmjVnYbSBqbHytcWXOwdZ5jjsEd1Uy/dxzngMDlIrH8toRwqP5M3kMAk
Rci+ufl1kzFil7t0WFvKXdwtmzwBboRXN0J/VPStrD0H4TTEVHTyRhiG1OlARKG82d5xqqEAiZHA
qmhGIowJqGWeENEgKPgx7+TsITISHU9kCH/R5kcyxtFYm51n1oH4fS+hy2tkt7LOYpkiR1MFOHxQ
AqXo8rSf/ewCBqoFnY7UFtMNvxnZTUZnaYD9qXCh7lHRB6yltQbeYtn7kA+z8qwGfpwi7hK3GrNf
vluNqUKkAaljvhMJTf3W5B8YQPx8ZAm26MmckCLYicayKZ6c0IoaDVsUpCDZ71R+U/T7GI8ZlQzO
PSl//oarqGVTUKywlE5zQD/idilmvKZHAV0JKdM1+XtFCuLFIY9JGY0ri7YU/a/hxyYOmeukehX/
H7brcL0xRSsPHdZHhmoRj9B5L+gret2/zgWQ6khzKl000unOwiufoSccksxJcKnhDdGkTxUHBCU2
NNma+9SthDtYmbYFl7hDRtSPxT6rleWbq259c92OS6nbOqZ3+UqR+vS4fyArvCYYbTF3wbxVBc6O
QNob4h/pxf5iLOO3rmei39Q3ZmoXbbNPxSFTDrVcfYuM0myDhmaCqVgCGnuC5tDkufVlbCURSs7L
INF6WOS249ExU0XgY0Rq0Nu5sENByZ0emFAtuVDTkgZVQfQB0QJHsxMrB71t+ni1Rckz3MmiyLOq
JIbLqLjJfn6+llaTnNKSBvIKz3b4BoJsRy+meVL2hKj+OLD1FTOaquRz/BS7h6ngFaa3Q8toGaSw
n9UWeinfoZJDY6Rk6Hrr3A75jzT6V5rMCzbtlxVfo+shnI6likQTtK2KcBUOE/6nxivzC9Js4N/3
l1k3rcse4g3C/1wtPDHs5ijSze1xOy0Pzroxj5S9Krx7PPiS/IBMwTq1rgiS22GkNWsyS/icF+a5
pj0g94Nrm/GwvbpDM8315uy18QVfWDlHsXV6z7vz4DEGRs58G4XBhh0A42A367Nrl45VNBl6RJ2h
HUA8sJaTSjfa31ycKto3nUDI2kN+c3D4Xb/ujXH3gB8Y7L7qeRH51cdMgCUmjCecbWAzq8Ewm+++
4WhE300Ow2DFUD8gv9iUXzv4KbiiETGihNhu6R89hmoRB/XNXvxaZLg1eyGWRUcomiD28OCOFQF9
K/iqKc4Pt6SlgctX4TU4k1T6737TJsdmlQeI8hHKLkDBxXFO2e/npwnsvxmN4NzQFYIs2pl7lX33
eSogss/0JmrAFPjjbXsWHXPLkkM+46f8NMtlYn0GwG9caNsi9zEUH/13DFVO3H+9gRBgdtdgaWRX
kbczRTtUO9Lf6loZPGbIyy7qBIPFCDpnsoXMsA1XfaSby9Weso8TyTbrANz+EJDcd6IvDSH0ThHw
fF2Hg48qKK7FCzktHbHrcOpmr49JDfH3zdR0WsmCxAWQtAF0x8PPpeL7yY3GzifUrhTpPlrXxeEz
OXe3g7uGnDj+ZOcKvS2+Q6hioCLR548cxmGK28CzIVRjO9M2D8GNWDiP54/5k/PVfiB7tbAXZfh0
hPsz0CqUMFTR11wBoptcZR4Zi/eq1nJYq2Jg4kuKBAwahuZHLT3vSMkXrIBLIJUsV7/wON7RnUmx
oaal+yF49az19lxzJx+pPQxIK1CtuE77Dpq2vTYJrqh5bt/m2XynmcqXUH+mn6G0gRo5oiR6WtpO
zksxzG7C9SAgtFxRKLp2Qw8Pi4/rQegtMouVFjDNmmPib2xeaececFOUXHsMVvcBxiTaVG0hERiZ
wcFqK01z3W9wxiP9GdQChZm0uSBoxryAEcXNjT/nxGK2KJPxO6E1Yn113//GhlX90LZS+YNVS2ix
X0HMOvYx83SzukxPk/UOWhBkmuQTTnelFN2ne7OgYJX/wQE1majElbnFqvhXheRvg+IYDNKaSjJZ
ufftEzfoe/jVMH6mjUAIVZEdm6TJDiOXwlCrxWicPwyWVnvCOcKs1bGcvnI5zfNvUz2KnNxe7Wbm
wLeAPIL5Cxx78qLEHvm/8VXRDawJG/jdhR+Tv71AP6TwAmADeNndqtCrVqmF8JJ/hyInw517uOBv
ujFmO/+Xy20OACSJlXLhW9JNJBn52hoT7tUNP2tiOIfZYE/2YP24G6DgA6Jui067xhFNOWaCqGQZ
Ci3ANa2OasT8QCPuv05NckAbA10OPI7FZ2fyB6YNUfNb818fqdF/BpcJ2qe8hthIJDkkggILAYGR
xRH7JT/p16EPiPwrq8SKW+pObr17yhrSU4BvpLbU/sAYJ3kqphRE3eQQPBkXD9C1gaVliZRG0bem
b/xRC7A8fE7FOJ9Tq2vxpr2sM/d9ZdlFchbht34x8KCHcSsTC17lf7PGtAsTsyioVHQJRz6LYdr7
j0P+RZ7mVNsXR9ChxhxGmr2X7LnwPmzesvUyPOxZntEl/s9/Sr69fHsXnHe33YBT7iUK7W23IJug
Q2i5f3LISF1uIhj7hFKaWmvCgJW6ad2WDE+h4s/3GWKkd/d8LMbt3DethMVOLdIO9kn3IYAtCSv4
04w=
`pragma protect end_protected
