`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jRtg+X5dHNhG7V9Lmi4i0WSBbCRXCGB6n/5KHwSAkL6C+EriJj0K611f2xiKT2Zq
bHmOIhvLh67rIDi5XoWuopn2bR0ikBWaIBTjgQV9nyO6Tgce4dH+g5h367KT9w2g
+40WLhkvzk4p8O8lCRbSyHpj5o5U5dDQiTWPyyBUZ1o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
sExs/sszj8zCkC4NuS2hffs0CV+U//D0vzqOzelK+N/l/QvkLAjJ5nhWf5vnUCCx
nObeck1Z2rfYDQ58eoequrNn21jm8WFz4xQGvH/3F4hCwaEA9aK+hy4CERRcoJJY
s5dumvB9NjW5FjUDwFhDJPDzjzuv3ayTglsnIFZ3M31LJrIRupz/jVestnKMQ/gX
oMbIv0NovI5YyjvvanlLR+U883iguToNVclL6pw5rC3fjwJ+/tbfShOjxXgF6wp3
0G6KO5Ee6PL+EHSyZ8thS8k9cbUE+urUudBjibTpmkqAo4ddOfe1ynqeEJy9o82r
C5jFPp568H8c8Wk5g/n0+fRgi0x2WWm7fIXX51rdm79h2bJ6hdum35pr+pZJiaRw
pbQQxf+2+4fBE9GYCokXSr51a+QGQWyLjQILcLYczko1iV6iOUXWyh4pXMqqreBL
fR2epJoYAm+6e6ZfSlWV8g2xhu+Fmg/YWu39uHUS2PKB1x5QpX0+LTRecnmmSPHD
Bn/rfIWrTq0KjxA8H6eHQc4mfs84Onx5M3kvcqmLJNRwJ5Vq2D4G6Q5xbnUrSvql
rFpgqdyqmtaXx3jsdGmd6xlejN9qU+JpqpCDwfz89MzlUNWV7uKt/NP3uw5Kwgiu
Gk9RrIylx4NayL3ntRo/xg/8VGs3F5tYi6jzck1mG+PW4k51AOjspQ7pN5TedX18
c1GgXgki1lw3+EYB3fcMmxeGUsvtLJllcOMCUb+6fkyzYCjKhY3cO+DH+Ct6K/v0
wWnrJ786Ygbp2SCNFhPALljFnMur/B2hLu9xkpzetERfeKeaqsBCU3DQo1uVkHfS
2nhl82oO6BL1066WBKEuNXwkkACmk5KEQbJRD2yBTYEa8KUM+9AXhArYC0x0QvUW
G1ZSHAaROYWGLZ9hb/SCGidrfGgHYaMVr6dZQNi6Ial62DJPUOo6UHB60ougzgAG
G0VWMYaSP0uu606uAjbNSMNyhQmNVEMKHsveX+Qxpup+AZkEk77fXLqYvmCKlwc+
AmKtGpwZuqkHaAEcoe7bsduezKfSHaHa4nvthBYsdHqhuwxj4wXBsTjYKj01Ft3/
Aoq94hH+pOFassb1CsdqPgS1I4068HRliD5WsAXKNkLzWilSU3a9e6Kc4mRrW+1A
JjY2VZ10RGr53FcCMgoYDzVKVeVNQa64y0Jk2ejz7ugOtrWgQTrTwOxigcSBfXCT
GMariV5ilRSQw94wRNlK/zzeqe1s576XxEWRuicSjmQctYhO2hhxiRkmSrT3NuLd
7L1Ux1o+Sn+p6I3PKo/BRDas5qARy8ZtwCkcVWh/jEmptQ0XwSKnLaDmWuC4Ngh6
aBGQNHmrDqKZe9A6I0Y7P9TQ0j/IQlWwQPTwcE91b9n6XjEBT0Lr+bLMgz5Wqyl9
WFQjuPY4J5GT65gBD34eLuLUBoftBfkBPH3yg5uCDyIbxqYySD7/2s0SDJN7oHoC
kNEW+aygoXwe2qV5a3dkQTvF1IMn40mVS3v4toaRhjE6BWnsIPlBXj0QCYp+H9qC
l11rNsw/sqewby+4LgconUVNWVFirRm9D6nHsQJylDXX/JiWxk7R+qImXp2jKsah
VhsY5hdqYmeckYAXVNmz7ufCGeY+JBEs0I8883lZ46V9+Zc0IXWljfnv8ELg/+rY
5cjnstl8qyhAD9ZJCr4d9SUQmrWSDQoUkntpBeZOebRG+ACh5xd0JhHku4KUFS4N
QD8cZRJiaTBIL1P9rYtpof1CoQGMpSalnD+gwJC5ZIUn1Qd6ILxrVhc7rMn/mu5H
nsH/bhqiJfpN3ufXni4xzooCnu/0ZkQXgh13GpHlZmsgCMBVPMxzqvePDIdCqGsp
XoByaj27AOSui7fxH95qp1bP5raFxZbJlWIFJsOPr0YRGa7Cz9DiIWzpf7sm3+C0
YYR0SwYwHJ/wMPQUozqpv0FH9hbrkt+UWiOoSndtFEl3AABzYNNuRugtvbyUoW9+
oKMTe7QdHFUadgTTIBjmtcd9RY2LdZqV0GK3TUTWcGuFAUETXdv/LolCeEFU+gD7
el2CjF8X6JjUEKgQV5BJG6PeBUgHeZDYLJQUrqoxMcxWIlgrWKWsO3HfwTXzfjaz
XNy4QNKCjcqX3KcOcLoMxk+Lhqz+gaFCa9J2vKusXwsJUhDuCxIaR20xKZi0pNZu
62hP8mEXS8BUdOWyKmcto5OD7FZV76p/IFU/XaQ0k0RXrmZ2d3rPnALgqS2o+R/B
cUd9FhEyqe72Rn68Uri5wO0/H9+ASyT9d56EjstTTmR9ixEX8guDFn+tHr9Kyt5l
oznC8NJJLevaeTVXj7IX0JQyrLt9fcOTds3WJfpek49od/k/4n1d9lkVT7v5HhzS
8vejNREdcEyKLt5ZsstTk3LBf21r2cnWKmlVb/83ighd6EiYppuYkdaoaPIu9lWu
d/IgT2WKlysHAnSk2YGJbaHvHf0TsmlIcpmSh+LFohBCuMYRYAwcPTqdx1TcUxk2
4yr55Vi0qQrhsXn8imRwKHNeFYhglExfJ4vTF80ygiq4szZGMMRIfLi1jMXd2pMZ
IXOlbhQ91lJhD0cvFsvSzPEJfcr1+JCYePfCH6sntUx3NCFmRmkPwSN/Ewsjgx5t
GHlRIG013iB50NrBmWCQjI6WNAFkctrbR4WFLmA97HgDFOocP/0UJ/FyZjtwcz1O
xox53Cz1mHDPS4AiXhQQmtML4O9OrnQY7/OONFhPpAoZAAgry/TWXfgG0yyO74MT
fTXN2AKuwlQVuBsw2PyAtjcYoLiwT5d9CMSd3i3MOIpZT0P318a1uSK6KdEaCeIJ
OHu68hJNyCAmTYc2SOlEt4lMCTeKdFktCGVNkzN+fM8ktFnMMNWSp6A4BCiBdghR
xvN97/KmOua2kwdTNA/fpR1xcECwYj6g8nSCfHwshcEUhPb9HP6bSdqeiCjxvgbh
s8xKfHnyVhCkou+WjFPklB39XwHz5L4uDmYcHLJXpJBPCEmKD1pKPYlZG/T5/idq
5hx/GHxC2bSPO22xlONTQ2ezBbJtDK5h2yQvNbzeXoUoAj9txZKfp6RuEj6xgQYy
DuyzLEEq+N+bYEp6h7vlVBAxRTdqQtFDlHT3B/OQmL+XH7tC2NMi6Lcvq0OrPOyy
d0yYXXI/q1H1azT2mcOxLZXM8Vt7PbQEPvfR+4jcAH/vYMXCm5qSPwq8Deqic+PN
qqpGMd4csqp+mnTp/yqu+brebi0MiUIpnOWZzaXuOxSLghMua2RrFIwYsSUf6QPh
2oezmYznEw0LlP+M/qSSxOibFse/uUhIgBqUlNsKTmjfzzSvI6v02Dw2RFY5G6g0
Ep7BVVK+YIVTAivSZ5QU/Ws045ECz/TmfoxP9dtBGJ9pUPGfhVWHRLl1h3FhP9u1
Cbnzhs6czBxDyoXXPTrrqmzYbYD+aJBxQw5CNpWVTbA5qVvc4uK9rI/LCHbZseK1
nN4yXedWKnVD6BQJwGjQFKQLOb8w/EEilWitVtsImwDZj9SOQnBb3OfCGqAR5Nm7
wvAplYnRBpqdcGkmZZR0wDftSB8mj972W2w3wOLkiEwKH3CnOgeAYr8XQGlNXE2K
KoE8H9EonqSgBdii0DxATMcbNgUEakkLZVy06LNw5c0L2x6nM52DET1WA8OEPmu8
kY3xW+wJp1go4vP9i/bMzo2NbpR52V4lokjvPhQZ3AuJZ8cJbG5QHBun2+5mpFCK
dXBLId1HEIF7FDsudVEHy6fiP3plNxAsojl4dPvHQCpEvwLUXR0iwaynPW3Zv+ys
+KxsZYM/h5aZnSuN/Vn7NmDhH3AIRjTy944nWbkh4a+JPUGSMEQywRvCWRVPAfFf
ceCjdZVUOLPBy/wDOm3vWYJ9uDQFPyKLyb14Tv80MvwLPAMKEJOpEf6rpkG21BxH
ShDi4V8mQy5TjFUdrjghTZ4L16Icyam1EFUQCmgmZZb0Oqi0Wk08yBi8NZ/S/et3
yXD7BfSWPePFEkrdNqHP4y0UEpdqfoYb/dGvUqxeja9+lNArNg0VH00XH7xK6O0G
ZgrXcQQ1OZrQNZKgXSpghY4vyUyEyexCoF+vvYVzDBgUb4/678jpQytaILV8WGWz
6JhUZJLKD/S3yDObV4ogfiISnZbXMlLWHjdvQW1JQmu5s9lztMbVSR15NX/2ajqM
4lTX9MIvC1VGztfkcJGBeTvdV2Bd8TM7Dg53NP9I1TVEUlQ1CY2HF7CCrXj/rzHW
f5Gh0/Dk3Dy27EdjbAyvecZc3ULJXw3WsZYngUW1XcTZsRoqsG1kc7RhwbnwlRjw
OyaAiAqz5qEDFUapB6GZHi6AyN6hQYCTCGyK2wsc5c++3Nbrsa6kb1WVLtgYQ30z
taYKmsCv9vBJ5kQB2GLnol8CrB8h2eGRMasTyVJg+J4AmONX/+spuQHfTMKUOAwI
TPsQMNYmYAdX/2UQ7Frn5fGrZuvA11i5ZFA5WTA98RwCkI5Nyd9TlNDVE87yraEg
3DV3Od4DJ4i4kPpPmWNHd5myNN9w5amsvTV+yPWhX26Zq9Kcgb1t5zdozdzVt1Ph
TnAuH2d0kNWJbDeEkPaDK3x+gZDq0OoYI+o0fwKX9htZZ+uoIir7wTiVvhGcmqbs
50o2KPrN4yWPSHt3vbbSi/wmnnxINlRaVRVZqzzm10BQxJvXyAMbBZdcO7Ti2imO
7s5xSMEIv/HSgOvJUpRsKaXn/tMrcZdYnwzNOeQ+1/GwsZDgqBHN+GB7INv/nSAY
CJ5PChgU8apMgnA9Izc6o7ibA4e3pxA52/uGZ6eHbhyfCde6UbBAqCBrjkE1gDGR
Y2DvoLoX4SJrWnAk5PiqxXjboSZR4WLkLMQpAzoCbyihYhuOIJs2UkEGj6RJhb9m
Kuleo1lvi51fteXZXT5ywbSlpi4zSfXAGmg3hOHEfQk3reV0YKpjdRrFFMRzTVwy
I9D2LOlLPK2dhT5I3uOFGpQNC8QG6hnMizZGf4duGlgM6YAya+RO3y8KAU1Q1R6l
vz/S9qnuJozuZexJv6Pq1XkTcb7BP3UN1z4GeQSafHmzhiVayWsIwbco8Ut451/Z
dSh2jkYvJ6qcTTYj0ZueRP1GfIfllORlIiEBdQqAQNFipclzINlW3H0Igo9yUj6f
9N/3GOxE6nWmLTTwv3qFN9b4+P9l4iguwl0DcYMWWJ+9CVwlZLRlq3ZKaAP/rOFa
zg7NPo7UMv+gVwoLX4ndtaWYSMGZvQ+BUTzsOkhaiE071JlczDHLsqoLHjAeV8Hl
8+q8yVtO+vss/p68fdvjYJSpD02uP7cz1bhvUs5FRvliwgwEpaf5SFORcTVsDed7
5WpJUdV2T2WJIaZAcnV/qALln1qf675uk8LPPiCxP+wqe4RIkxHn+XJeiDwyL981
DW7nEORMiprVVTB1k65ely5bLB4z8BZOO3i/ByJ2uf5H4itwJhFI+hlcnT6Txy0O
lNEF4jscrj8JKTLSuKt6TzjE6SMD/UydiDz6l3bgur/Zr66u/y7xRYF/aeQc8yov
aAiATBEsvejwROMYIw3HgScsoWsSbtklfHcanOJwDDvWy3n1kHuNhOt8vQCMQia8
wpKhCu+esOvD/QNNkqIxu2e3/Fjy/mQTnH8MKsbp4h1dhryNvM83B+6O0GHZNzRu
5ZKh8VON6nqHW7QUclIJR/7VsjHb6/jVRnH4wkPCmmbvnzYxJA/AppK7rXCKJFK2
Z1pEOHgR+W6OU2MWQEn3OhykgWkDF/grHQXeXXyfvQUAiG9JTqh58wQAXMlsxnmR
EOcd9KO+URYa/TA1aTrTpol7416OKvHoMM078OAtcCb2xBQZzOJkQwK3YZY+DGkM
qfY6fDbyyL9kkeo9gnauUrcFdoz2VU9lTDcSsaQKWlcs8xD85zbsnDU8oHCWliCi
gE7vlXwTw28R/FRDV1mSW4FBE6GNSyhH/Yrl1nr4iAcWYhtGi5r8rP/VehSz04xo
Wr170nCGOVdGAzuJmUyQVoMBGfMcJVKDCmB1jIx5vUWnest3Y+X4G0ctwVrH4oim
HcMS/xOrtR+XBTZ7pX6BJ5ODsJQ/t8JZkHpqjTsh+CZFndg0WHigWj0atlhOTsyS
SIgiAaxptgg2s3bHaYmD3CNVZICXDipVO6eamescQcf3Fz727uqhENzuFNLkZTuz
IrrA4/C07Ud3jp9Yoyb6ya26KGSEwoEErjNiW2f8HkyqBJWI3AHwt5vDuy6SVF/c
cP2hCBz/OPu8KMMm4UQfzLFVzGzPttWCvBaq4gk63lP2VJNClQelWQvkumfkG90/
6KWMX7o8F1hPk4/OyzNFORuwVe7zE5d/uR/iY+JWOdx5mw//qIWWOvOQcjhfeusw
ZiYg0OXW44V7DCcMpQakKUbRv9Bn94c4ImkZSF6Ecteu/4LVUNfBaJ8/xFIkTodA
NBPZpnlYmCQdDbDDCKF95m2YL2PO7ajprXobHNJRwYcZHVVv2xGqXCtgjK/ts/Gf
WMhhbDNxjgyUP4WQiOcmMV5zQHYy/aWTevvubyV3dFwyYddhDtvzN2S530I1rKsj
BXToQPUbNK/oFvz42zFeeHclAGnh+HKmC9WiEx3TYwr5w3uLSZOUG0pZznsJTSC2
Hk4udUEhjBPU7lhAWMcYSpijdtXqAFpNTISoMqlpsMDU6FfLAYNR7HS42OGZe2Au
6LZyOsv71pRzlSssCF2Bh+JgctRJ/CfMEWICuVZFNaFWOkDs4ww/awCqyYR/brjy
AYxpa8rUTl+dG7f5eQgyQdW54QyoPGfdRKNvhp7E+h9d86I2HdvzqsnkHdIswQo0
cQr73zEQRFd7dG/jATpQGPvx2sjlJlEQ9OGfwfwW4FBkgTBDyS+WaHdY33QsAODa
7iWrZ/TxrFuiWFnPy0wGXspXM7ftcl/DbjwgzZR0sp9oc6gRXboeiadQyPjFSHzV
aeUhbKJBFYIH/9NBvZ65vYiaMdTlHlONjdbDu1lBU0dfqo2YtG8/y07AbtcX6+s3
9oWvcyc/07Dcq/eZ+P1Rn+qWbf0bmdxzVHpdsQ04w0HGmLt4cV+QWudy2aRXNF+F
+qtZ1sA+R0HXK/a3YBSXalwo4XbW1LkCrDYJWB+BCwhL/07rJlzXLPQvbZvTYiI/
BWU3jxOUXomcgbdMlSWYkxNu9isIoE7n/dXxBROhKxcTcEziroSU12tfRhSZEsu9
U2BXfZFa2CuN9vcPoy4ZJ6Kfqevl0jRhh6dW8JNjXppN5lx5bScSCl93VEc99AxY
hfQxwxXmBE7Ccc0/k0dttMRppI8i3AnXkkFegYka6wTIazU1Y/+SxYXBVl1lEOK/
Bej1qferD5jmGZ6HbGUaX55jZjZ3xCLjTED0p16zNouzFTGtwaxkMFtmx9iCxiE9
1jA+AJTRxgF6buRumyiJRmkq7iv/IAF2MfuMmXYgKoleXFLzeu4WnHf4n73r/jhH
lb1fqcXWemhT3otJnsl/qOq2Q0LrWgvY6ttAzLrrja1KkfzliwxuYb+AIGBRzxYL
1diLg03xBKRLy8mk0wUuoK331LzpK2hVg8N4wnSD1VUonEm82/YWtRT0cE1lAiWC
3NuIhOc4gt+3t2sNlptBsp/c4H7grL/fLPS2aIHx23U4HoY8Ehf9PnZDiuog+7qs
NEoWZvgg2BwoPPDaBf3dFtGQZl+Ka3FuGl54WGBWInmOlpWO7MOot79uPgHJ36BY
t7VMIoJPtjRgb0udwHs9qatZgakA8TF3MVFLUGmIcR5xeDfcOLyG69DNvmjilWac
dydWE92AxuL0NIpY6sdE2vORKKx0EbjkI3q08E0LQ2Tamxcx14qoLT+CHe4JXp7o
JjB+mzvTgMlhZ2ufDkv11AZham8K+HUCOc30ZOzfdnKFJR0NLFtkTl9fZeoDljkm
8lMm0lBgNkdv7svHVBvdG8g4o39kWFdeZAfdMWZvPVH+IGCNqZ5sf3OSZL74+Sh+
9Y4StbrqBGJqp7WY/tbtxzW9BnswL1enI6T8wXL/JpCSJOOXT229wnOyQGOtuIhF
dmHAZpVQj9FJQYO1TQgE2n1M804Kl5K0SKfRlSxf8kQZ9MuIrY7E9wFEkZ97nPhM
Bnr/jz5HOrkcAW6kRVKMUc0ck+HyyqX7DPk7TXPGcQczfYtXAfJA6RZBgw0TLBG7
f8sA2MghaFxH1nJYBnjaTj1ay3WaapC3uIWaShAAYbmytDmv6NlWeJ9iBOEL8QM+
fssq+zh3ndAMXVFML6FIGM+rOzPaNV3ZvanjUMuUUTM4FhSLxkI4sS/+Y8bznAnl
JmuAcORwpHiJNWolhOzbUgKlV9HPlZUYjZ8gQU38ki2eFomakHavliYFQOdeo94J
1xGd3LtowpDZujp///zOsph46wfAnmUnZaCj7GEmIVKBOtoxHGWobYYmOPpDcAxo
UDc70q9sLLIJcs6dKj3OcmodKWr3PMGmheU9CkXtdFSPT66w0JtWLmVXNcDFxhws
WbcY0qz60pADJDufTQCfJVG0pCc0aPpQs0Xo8iPCmTMs3gVMcsaCPCvHmJz3iaeH
SXAiPjRC1SzxIgolJNjaXmS7ufWUfAxzm9AGatOIe/r86Gp1/vpRwFo1eaDLZrKa
KhSaf0CClx95ipQBtPnUj5YsHKgcStYLVa4W5rFdSld7JMYXXFcS0sQ9XsvY3uWF
jzmhdMdmvnK0qRMXd/oHJUD2CC+ClyEBoNINlzhf26BJpNqmBBi/U1jhxLektf9L
iA90czmi9OmgYv6nelg42KbO2prYoOKQpn8TpnYXLEGghtC2fNYiOvhsM/tzEpWK
zYVlWUkdrb/DxJu6SnOEJXKeX30Cp/yAjmg4Q6UKPzZ5/A6o5WCJNRcz/VZP2aw3
HAVJBXzteMnBLpi1N/c8KhXmz+7TIW7foRoQKvumvYErvuEJRA5n7DNlnUTDGVe3
c8Np9+NpPdSgxM0diHxwNThfp/ho6EhQmI7F9GL8h+eBlsGMM5hwrOkjXQVHY0N9
3TYlHrqOhK4bHxiecoRuniXOV3QERFnqCWVd+gIpfeNCbIzGy+/DWzU7E4LrOlIW
MIi6ypBO8w8DmvKtjOk0EXJL1RNBKIk5LyNZKEFFZek9+3yY9xs2o960Y1Lm2+Fh
JLxtZhUSgzBrkiq53hoYl+zmbSsMeY3DKmmOydFIvD/h5Xj2xpf3Ju2U1Zlz+SfT
dz+rKv1OWi/hLmw5Ei7nL/TFxww5pxdaoIuM7Tw/1lr0MMgvaiSg5av/ZTUD8nYq
B0OgU6bq+SeGoFIE8wy711ccmm5lqQ0OaVO3cAo1JyAp1wEnLBg/D0UU9J2Y28Nd
oFloO6XMD5vTlZWB6YRfPDOfybaG6WJG7N6c2UQhjLtvLxyHrRsPUoksji3TnP91
UagZv93Frw/CBeMIi7DpTej6wOhmd/KKJMMBEu4A+0HftlQzpjN7mz2YKurOLYfB
ZSiuGHyKW3zX5QwZtxCumE2wyhA7n/theb1TDeW6SSRLa8wYxggZOsdeN/uSkQyV
8wEop0CzpW13nH9teLern5BlDIG1NvdsdFmpw9CmsWwZsFe+ah+N6sWXYIZwSB75
bx1TFllC8owiVBSJuhFAEfU+qEUQwaBfj3JMJwe1xC/c+Gu4yzJaTDr9JZALwykv
1WpPnF4ak+R7OmLjmtqSJp+yoJlBjM7BOpNZZ00HKj4SnJQ25geUtJCbUdyXsZNb
IxzKYg0y57TJiS8+yNwXLBD/dv03utazJk/lcieBFJ9mu6cYv6Cq2nlpBcwed0FF
vPCX1igIUR6gyEMGV4aUhWT95Urh/TldQq7/wUdWC/SH9pe4krwinQ81oK7kTa2C
1KBd3cePzfbakA3aXQzTh4JmqoWwoFpfROPnpuS65i5Ny0hccikTBLB52kElWTyx
ykpboUh+fm2V5Nz81fHebusbtTLrNAa0pyk6DiALG/4u/rZ/gyAjzTKfYEqmTOuM
I/2tNp3v9/BON4XUqibTkLd3z7mDUc4paod7pPOkGz4TqXROFvMLlE/ru4RckS4s
Ak269oGWUuZsckTVFSKlN3yJRGMopqMYKzJwZ2Uy7F+jZFvSwcgU0BWck0LivqFE
HAQYF/9c4YOGB5F5JYRkgYzw+KsZlMIdoDx6ZBft5bk/Fn1xtW2Yq2dWHSKOwaIw
6WoUeioSJPWoLkhWjNSHfjUFa4Mia3msiOqWhPs0TCVKUURwdfWacP6JH6s8FvEy
sBXxEO+6ybgWTu/FbiyEuQgAGAEWMNDakYYuJuP6LjisDuEFwz9ck20e81spYG8p
pdw/oUHA/9S1Qn70lEhbzILnj74b0A6jOml4RjGQbAdIV/ppif1I8PPj86hth6OW
UFRpSgKJbTydCwxySWvc9cpTvwvmYNaxHi5GihRHGZGGFBkT9GrIL/zSorZ2Zb4K
mzzSv1LLrfuWoeiLuwPhzxw72jFjG6uvfAu/cyoJUd/QezczDIlyNkY+fSOf/j3W
4v1eMsgytf3OL1iSFyPmeFaf2ndkMyzbXjR76wkvTnibuwMTYGb8Mw9+KXBaVRFT
XHx1Px1PucyEcbUDcmXHCkEKLbjGSIfkAtk/2GaRwjah1rKLSsks7DCMja7/kY1o
OGSwJd5lG0j947JfvEOy2HPqjd08czchIv5h2Li85OTMyNVvat2cvJP5rmXfZLSI
QR2d/7coXQsqo9jHxjI9oON8fSAux67+zWiBCqM+NphhCNY6D6sAje+aehDCAREw
0NxgCpbmW08K/9l9oAJucGyqsYctaw2OkZR5JoQzRYIeEV3bEUsyPAm16wbX5meS
9rzbisgCPe33s62rkZtitbf0/9ooCUaYU8oxJPkv4zlSLQcfuI7FEqk3oMzrSAQJ
qEzQIN8/0Ox7mtsdVSwUm8E2szAwoLnkBmvBUV4YV4ygPl2mCZvlzw0gxOYgjsGq
N1Na7PBfZZ8GS6u+V/nBOFG06BTkt3sOqGYzyTfAHxSQn4xF2G/huweg2Gm8CHD3
pKpJIqZ5KdJHlbDh10skg1PgfYbbrqVmkn4caIWzmC0798G5imFlkhcQmoXh+3uI
e9UfuT1rbLv0ZxQkUKF5nsRcD7fzn6GkBXIfpoF+lvDyT3zYEULD5VtrPG1K4jG+
IY8uQeQD0hNY632m3G2/Vm0Tw9CzjHzBOyW8X+xFNMk7zh8M+/+niKIqwl47ZwBf
3/sBPqCHxfhOSY1AVJJytEVVnyZbAti0yzC7GRH6G/UpivHB/1duP0Wfrg6ovxfE
tUYNVCB2IoJbsLLaYKnLxD9fW6bESvaaFGm/84m8Gd8QAW2q7KlAWtDG20WzjTGb
oUvD6etc9YKASNBr3snFVd1/klcrzbIndeuS8d7wUhsWlW4qQcZjd7vGZV93szcX
zepe0/DiMFhnnvNGdPklDMP8stLV/GDHa1PoDytKeDqJTs7wS4NNBSdA2RYG4jPC
xYCRYbE4VogYjRIW1wLMcCoEcoG63HqC1zn+CziQlGiywRPrqpRejdLsut8XW8Tl
w2up5G0gkB+7hQxRHSLJ3Gr0mEhCjnu3r0yITTj03sIPd2ebtW97djOr38td9I8k
07UO8V+JeEzJgzVVQPtNlV+O2Dzg957e1/BInnuDHveg6axiryvsKgm/ZiiGnxct
rAgLWYpu4kA+B80j4UT0dsqPypXt1TqLJAgIC+4330xXzQ9ysUowarmJ3J+V64SW
qWfsBc0j8qx6OU8ACz1mtZo1TdeyFrRWnkXxyoDNDEicbvTj7tpBt9J2eD7wQOnq
bwYQLz53ThLSsbjXqEiX65oNu5Jr9jXErEWMmAoXlA0uDUNdwE8ZYiL40jnMuiiN
S7kDHsr9scGf2tkebazsdFkvRltv0YToRS+awwCWQSRrjvSEQXYoSsIZQgxE5Jul
86s9X0zRS2NMBi0bfG+Mv0e9q2Z2FekHrvn3n/uxa/YKDTg7j6MJw173UOiD4QMY
QF21QDO7AFlUup2CQOApBvEtkyz/BcjPmL05fKi/+6I07hdB9GkbZyxGkPROSyYY
M5EmK/Dl1jRHlD53W6TyHfhnX//4b7E9Nyfj+GpDX4nqn9KwznHxFzpD+wI0O2xo
FGPELaJkOCvbuQqbpWMXEQ==
`pragma protect end_protected
