// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qRBd2D+3UBmc+BJ9fJwe5hXuQcqyv1sxKRgQN095VxcGtQylV//0Ov+Mq294cUCZQCId+YZ68HqB
YvbPLLbrhUc9up3WxEqr0ctlX8wBJLJcCRMe8TOS80dCsRLmh3J81X9SY1+xIcr0GGfVJ1zOMT+N
lZkR0geJaN6v/0odANt4XwaoxgLnoD+kggehGfZrIgp8tW3vaVG9J3MCaVABBQuyWgEfJz9EOz4e
Uc+iPsUBCfaG5jn0kCY4OQOSwaglSCYmbmicNm4vKA0Nsj9ESdA3JBhEKKTcJ/v4Ec/Gy+tTLVHY
nVrKjFykY/dskzwMnQ5oQbtmsmyzqzxgg115mQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9936)
HZyBTouxAxQffVZcUqB/QGCblKYXRAUPJI+Vqjfd8h8HCUyw6NMZzGzNU7+4B8NTitiOyWAet8wA
Cxx4Y3VGCKt4y2Qe/n7guSSe3IJKgNh1AWYRSurIJlDsAFI7A+qd6V1o4n7MIdJCuWodTkyLFadG
339zY20EraOn/lgOg+ZVrzNk/Y5d0iHZsppDKWT5/x5fOFU2CkwGtA4qzXxLE9jJEVt0CYCFtuN8
4genhp00tU8I6Oscsz8sX3iBQt9NZ1q/JZRJXwUWs0nEj2IUcTcy2SP+hyz/ypI4xG6+vXeq/yuC
5ZH5lYGfyJ7RaypdDOrjk10+PCwzpw/C6qn0mNJ/Oouj3g5y5m/NSVN3CNrgCM9+sWfUN7ytZmHd
W75I/bPtNaojOwBO6ZTydYvVVUPnH6R/Tb0g15Ti9a8qVdf17BrQOBzgl84CuQPAwRq5TNDQfzB/
uNQ4EZJ1QtMpSbkGfnPMiujdzjIGUP3GA1rekDTayWFL2fF2BPB9738JzNfICvqmi87xsxM6htsy
MSlYYRR2AWCUxp57m8df5zLTUhhExtkI5PGZvyGpqftWOHujwQwifgtzzEa+XSL0/K1nd3k0nJ2D
BpnpkRNU/XxSap/9eeDaUEN96N/EqFXetAKVLqLnw18NvumMFWbqERnotjXvc1ZnSSB3Ju7sndPJ
M8PZ/vaXVq98UIndsplbz3mK/voNuBtmwIePtItXCz52hWIWo5VZ7Y15ZjxrIQVNoQEpYgQKk8h7
EOIHbWi5dG2uT4fjlfu9ovGvfjiVDTfnAtBTBrACKAjitoc/jPfW5z9HAoUOMP0vxODD3XKVRCdC
UIGkQdEeUbTUuLt10YyOgUmAp/TQuO2XFn0E/Y4dLD+86p8zGPB/Wl+uJlG5S1+zv+8TmM6/kN60
wmIAp1XM74BZUSNEGjPWig1rQ8bnMTeOlwRZTg+VOPus6pfDjLkCMr8qE1bMQYaTlzDIwvwCfNks
4d7L8raH/7J191KcVehRp1o6pfRil5MyjKfXeLjR7tXtCnfO24GhTPKNnDUnOAnva0MNJrsLPlWl
KIYgewwdwUa5zTwNUiW+h9phDY0BNXgrHMUlvFExhkDh+LxMHy3P+ufnJN2+CQnYJev0tdXr9Xl3
1mweu+88qSOAJcHHOhB3KfvSWE5EavjWUwqMAwWtNkosifM5xB3tEKOKk2xv205gnZpmBnhRUrka
ICzipWzfCoc8Ohzl1WmK88ZKdtu77CLyTXeQA4JKRSD2OlAbVWQp/XIhlEBNFlQHFWFuZeu2dC+/
MA8zciSgUD2gIEvBgs2PqbBVz2oJZKM+cwRGdpNIn8rPOfIqTo1Av1ij9LAGpCpxuHgOF9caWlRS
ZgoaURA1PUTPBQPbYW6Xg+P+sOjqAJkXB9C5tn5PQEMW3TQhM7CjI0vgGit0ytH2ZGFZVfmSGHV8
XJIlbd5i0tMOGcH0xikPsKQGC6kdRwX7LUP9zGiXnSgwYlCrGU0T6P6Se5Yt8wnwxNA7UfKRZg7s
iISR9CoFvpfddX1uTaKFr+pqSx9ypWA/4DkwdfWpPCAGM/tybtQ3WsXxyxd02B9bLATyfbvRiknl
6Ssoc1Wf7RoNAEDoxKBSQ5PsKAV5kCrT9iBwAgizd9SQT55Ll0VQxbxLMVzlzF8B1GpneBs7cM8w
9Cq67tM7H+grXqRA4Qq3fdMxuTgfrBiNRpSi5s+dZZqD73HWRPoJE6O2IezWdqvPUHTmLFZLmsRi
ksptCkt4T0eKgsQ62XdP070YFmFGmopoBYlMmu4mY2WnFMy5+dM2FxjJ+4CHWPHA5gznU3HySZhR
1E1I2yjfy8TRV5IqZ36XOeKHlLuilWtYol+tRPtY/uwGN7gsECY0ztjduXs3bkCfoVXBnt0ur7T5
dmNBGXmnwsCQGX7WEfr/4HIHJr5Sp/MQkr9+6I7VaNjQVS1AKG0K3H/+zj+NFAmOrehDNmRP08jv
IfgvXGAhLDE1VbIMEUq/z7erA1obwlg8KHWpSwfuH3N5DJh6r23DMwCn2ViGGPpIDhJ9Bdgt/VTb
JsMUMnl0Vd6fI7IwLIxh+qyCjKh8ARCk/MWRKAEL5CecAhzKGBCNqDx8LW9OSPD1MHyxiolrGDvN
JXgXh9PoeDF66DIwmqkXLClQijOaMLNhyw1TPv/baeZFHyFRcGd6IXYZ9CmoRnBhSFewm5q9ak2E
LNODJkWESEl7JLYf5wnzchrDV5C2DakHwTW2D0z6vwlBEWtlsAETtRLkWiNn9WIUL9dFP5mvhPUm
W4c0SPdTIQMK0tqwABmP1vLSmQpnuL78fkpxhK+DQG3lHc7i/layyrXY8L9cQE0CMZpFI+GR8nTS
+xFfxLYtJy7cJ9r3sUjFV7SW+TuzzUJ4C1dDNVbPsLPXFeayDqWDNPOcEA8UHo6imac6iwFQZE4E
kAUSIEBcSAR6Mt3je7nlLuk2icdlB8mFePcPYT8x6NHcjfV1RgUBHjOrHUGVH5dXVL5A4LjQqcBP
uNIpTJ++O+0XXFpp/sm+o8iveiK+q35qMDAxGwzoPgm7pr3goASVQ7VrqonuQT+CILwnARJybZCD
RjbB+krPM4hw6hlvKIxDRaV5mZeXZpHPpc/mxEIMrJmDpVVsVDqK0zoAK4mU3KQJfQBsRlDOD3pn
Ro1c3VnKgzWNb09oEGm01sW6+9KfwT5hfrolyCcyw809XaG8QpE7ZVqMmdAYrvQWFH91EoRemVqu
frlZjLZJIRrFLmjUQIVmCgLyngYuqdpB7WQ1ETofb1OmBzVImMHxMWK7dvHuc5kUdrXp9JthKLS7
Vd1bazdMu11rXCLYsbc+Mcgh48myjYrL/D7US/zD/7uj866AQFil9Uo+ENkhk+cCahJ2a7fJow9b
eWT3doVKu/rpqzijwpAP947q6x2NadGusH4RgWaN4syuH3ROndXqDgCgbpmeeY7DyRBvk7E091TJ
Wj8td8UtH7MYn9hYJeEEvb08u3VOaER3uZNut/XZ+ghIqAqqyMwzXIhJTV838XU/eTrstGVLuE1G
r873cAJwNnJDaq1pzvo9MDLtsXKctfPvZRMvTeFFiHng5ynphZCxRdP367kDceo5y6uaGLH7Tz6j
QNyTp2DYDXOshLuURvjnim/DynAWjas+sFlDhkXhn0uKEfMt4IEmnPEBBc/ZHMw/DexFEU2NsnnS
tYT6xv6ZE+EA8EMwc3VHmS/oQfdHNcOlXAMMnyg3W1wAbnVKIwXJdiYrXS61qL2dhi6GA1Lnc6iz
coJIPW/L1Yoe6SDGbSeSzpfddiHoAyS5kqWXxP4CMuOptf97evS8OhMx/DqeW1mmzqNZ6mJ2Hh19
77IMasFeopMS7lgejrLsLyLh+B0wOgEHLV3hQTlPn1/21RXrgmzYj4H8y1Qut7hjGCfpUgj6qNCF
A1VF+QKEmhJCk0pIEl46hVsont32ZpHDLoMrfTQBkWR6+pJVZMbF88KxyWFpAcXoRT8i71/AA57D
keAPMclIg2rX1/AV9AlXmv9Ge1pa4GqxvVlGP0SCLTXHCES/xx8ECXfnWjYa4n4jdr1D89iWRB0v
v12OAaWgiGb7rjj5Ofkc4zlm/HnO6gBPC8yJL8fQLZoM53cd0iaJGyHtSS7Iu9qhdAC5UhY+l03b
48qQGdycxV6ucBoLb03hS+Dv3Ay2Jy1Q7IsGGXfDC1OwEUAPLSI19w43njaX3NdB+f71G1K0fH2n
5O1/W3mog4Q3fdKZsyI7BQT2J/kMao/TEpDgTAXbg4SglqxyDWcMcN5dj+784O5sXspLI4Z6xwEv
L+zPsl6Q+q4M3Z0qQTYI2YwYK6dc8nVTL4yvHpjUZRyIjYYBHivwU5WK13Hm1a6jL2FzwLfPr+sR
k6uvMbQrKipd3mnNO8kMLYhUNiJRZRHpK65XbRSXS3OgSptByq1IkLnU567ah+J3Km6dwEuWpD+q
5vdTyvL38ZYRmjGuuVFYOPJLC7AlTMtSk6GSdRo9OuvX6UcNh6ICra79XyHJhN+TvCzW9uOqtXLA
xlpjAEZH07TlOdzyN0UrTkpheIN0OnuEqEQ6tRSMItSKZl4hoxgUS1Ed4dpGo5S1JfOUoH2WL/OG
l1RE/CV091fNlD46C774vpDF8wRA0z1ysFYH/9hC6qqSKpfN9FO9EKpy6ekL+4uDJMzeZqcBpWNv
4yd//xq8vsU6hQG5GyDJE89MdoRunTaia5mYoC/A1ZqX7ZqmKpVJ+KZAHwzuuKxDhN4ATfKzN4N4
mYyx32fPRby+hMZGMz329168dH526PRcwlJWew03YU/zhJt1qp+wqFaxzYqxL0RBNzmUjV9YyAQc
+c2/DHQhFBJWCQ3xrhkKg3ZIO3S1QKNAslh5kq9PYFF2GG6KnM41fbdxyBwH82GZTrcv7kvXZ1MQ
C+nfMNsqfI5u2p5Mn+Eoa/GKQuTuMZ5aXyQmDlm/6N9YpLAQ3Zx9cXixRtHrVrne/Zn4CPnv1Enf
ADvqK/7bDf9yG9idMkwQLCBmp07rr7ZnPod3+pS40Eo/eYlVXHNl9yjhIdk5N1ZXNW724icc0f79
ZEFXTKI85pDQntgi7HgZzYRk1NVOULrF4qMsrjwGZKqs0BLKY48T+tcV/GBT8QMOiA+wMuIadak7
b49SjiZL8VtL50TbqogjqAH3OuIG6qufkPlTKWj+TiU7K4/t7WgiuOe9j16vBPjjosa8EbulfEOV
dhqVC8eUzxlrA60H33ynKcTws1YE6SSAIOquGOg3+l/9lxWW35wrVLonHDaOfx0Skga31EZV2Dbp
/Zs2MYrdFWggX5q0qZiz3Gw37rL7qjcTsgkMz277PCFd86MqFCgG+EXokhfWj4WfR1ubX8hi16Uc
1/3PZTbrAIAH4PZXsU4qDcSIjOzXe4jI5sFMLxK1lwl1Q/zaoTrbDYzA1k7l7lx4uHHZRnOLS0gc
CWbRjn6sHtueed7rrMK1qFqcsQS6cIgqGgH0FxjTsgKKRnTjltJMl7Czwsg4dFQTanZj9aaTebZT
zPM2kuIR+dh0h8/KthbvKCA2AcdUJWymjkUoS8PI8W3DJZOHhF0vH63l7CB7u+ne2g2FuuDCqCBY
qgQ307Fcji63GkWmbwu6NAG1UXx95B6xl35qaAO9SI/8+GuUC3nx/vWpUlnk7TGAKHCkWBrzrf3I
pHLMExn3VpuoORVzo22MLRzhjwegM6qgdArXl2ruH8mR7l+16UF2yjY/OOAVYlkevX9KtIAhG5gx
VILSISzULSqirQfjB0DqjHGXIN9HXQAx+XOobl2wbMVx8ATj+Fm99CtEIBaAlsZW9D9nLry3wTU8
whEBlWKgDFeTu93EWl5jrW4MD4U23J2xIalIBmx5DUMWb4IjnusvvJkrr4tmPTlith2OjR1X/ViH
L3fh5k1XAhAdI5Fi1F980QZUvagnaROSWN6+Lhn+V9m0W00LtXbuzLkgUImZtph0vm3hJ1TA1cbg
0iMnr0GRKerZwq4h/35JbU5+Olw4Wz7FKMy2lF7I/FXhFNpT8NvNsQhyIhMwBiDlJIZaElhTW6bT
B0FUdoj96iSn7jWZYr16RDBuo1rGMkzm6FwgzwRLhUnUNXS470s51CAwFwDpyLJ6wnBwd1BSTLwR
fx05rpD+pxhPiGr0/WmnwhtCcOJMsSx/jsb/Fxyz7hRxuM5RdQhuNRJvIQwykBHuRlUYZwsP52hj
2LkeufSR2OQDaVSRCwqIJLBkp04aufycihOjnZN1Da50FWi/HZdWogCM1nHiKo7YFRouMjHH62D/
QQlZmK8TttZxozC1kXl098O5Cd3plach/U46k1/KL1A06GaynFAxFdKnjmT7GE4zNgS7riRm0S5j
Gj9uULZGtVgJ9xeASiyrEy9F2W+muu33gDmMKzorO5TIk56pRdMC9e8OmvDGinpoR0HChgMA98IN
urX+WIGEMQKyPOaIUq2q9DwXDqsnH3oAblkRb5paHnUB6RyLjDHyB8ks6pXVrwyqTUEcTUcrIstp
lgRFhExdAjiapV1xB3A7qpJ+Q7gmrI/qphia+HZWg+a2L6+oUkuFH4a2sjWegon3pxHRxKebrdzL
mtetFSpMRS/NAfeZJrtFCuuu1+PkAgz+HDgnuSW52cGXEUT6ATGbjVms+GObrYdIA7U9zwlgEyHZ
CTSpIX8re/Y1pnZzP6KeWdZnf2dmg3NSwCRcMrBLkxE/CsTPBLHLLPnu+vRZ59qaSo8Loy/CAF9R
APYmXKCen9vzRTamQB0lvT0cRo95F+XbtnVLjJ6uOfTmYHXcRInfDHYC8Sgp/N7EeCmOvV5rYdHC
4g0wsf7YDyhpO3pr6NLI7+G0DBtejaXVypOMPz5GKUy9UTCi7Z8AfkrAd4upzid15RnpfWpxcXQo
wNBR6hsSI5m5ttOMT8JF5ETpFF3UxOcVh57tDDbkLYscBoW1z2ccKxFnCTbsHd3/aDgNLLHMS8bA
fL77HKBVT3OYIA7CgYL84W/1n1T4KcGH5aA2S62ZLAncS3M9Q4YgM7gzzzM48K1nIKJjXvOjNdHw
frwZFKu3L5lPCTCY8BOj+vqJbSASJOkdb9D6z10nEXB1j84utAyFpJfpW9gieS8u2EsWTo0iSUvi
/5rH9RujJr86MXstday3yz+ObEoIXTe2XhyyCeW87hGumLIP0AxFvb5kguf50KB3534F3TSxIiSA
5tWA9Ho1zfX07U8r840F7iGY4KBc5YGVnSO0FZvhT9IqqiVnT6lAK+mN41Ko4vVAxd2WH2nPrGE1
Qyn8eStKI5wrAiy8hGAcLosrBMypqRH9+PcsxoyMtl2+9UWik57HQgfAh+YM5sV3BsiMT6C1Wg2h
t1gU+eMCpO4mB+rDtrXyvaDISYTtz+5u3OyAnKk5qQu/ZPN1fsr+Pk0a5cjIXAKz09gNSqKI0PTI
mEXeE4ztLliPa2iImS8Z5P59gz1MrkUp/qkO+i5WyifRs6GzrJ/OpFUmUdUC8awfQUe9PQX1yq8L
c1L+sgq7RJXX75z+BT44cE6BhsJGCDn7yUn7Cnc8TBpA8xYW/khFljf2NncTEAjLrGvCtAGLpQR2
H/ujq0+jmbnIth0OrRcNNi8X6Zdnf3rPaZLedc28yk8rLjkw53rim2o2XkAuUOb1RoUWz2O7IcQe
bhNWU6F1QdiiTeDQnHhhZayQtUJ1wrjriLe1I/Wr94TD8oQcgtwaQLQJCph16YRM9MfEpvmUI3Qx
qnTogJZHzQ4gU0bz5EqD1/JfbySsq7YNqknjJGyafJZj+GeySTfpcfS+BD7cJaHBTC0bxQhL+nG1
qyXcR7ntY0skZ1+Adtzjwaf54uWhIZu78rYCxlLdtmGEsmyRPnkf36u5922d5ZdJLuHeSgd0evdK
t5SVcrrwY7p/tvJXoU7nkGiL13X7TJa4KM5ZuAs//8h09oLIXGyK9BCPx7ornwY0zpp2AK8Gz04n
OY+IDNhk7qpBKGkAfQLT/yEkVAJSi/hnowXCAl71h5vUOcxixJ/Oi+80u0HLVFmsKmiKz3w5UGPf
E2LXk/nO7EAIPZy6XvRSS/L+nFqzgstSoHBn2KTn/5wBFHZlVh+VLHg8Mcn3gqX9F8D2hNDy2s0D
bSjmQocWtSdCXFbGkzumvdHvqkxs06enTvqVH074iHltAHN93n2wHYt3WiENECd/d7QbKkGSLI+s
7ae97lOFbRWVBmdhqggJt4vJQ8ofn4n+la0rM8bkISFn8NejuAB5v6jiaoW7VCSLVnLYg0nuQyKs
SrFHcUDDwTrD95+RJSzxS9XPmIcCXsVsBDgq09UuvtWBIbNs5XTe4Oc44rshNkAmR46I5ny2MDCZ
/yiZp50iMO7Q+4XYMFo1JiG5LjpY3p4r1M9G10KWH0BZLjJDnzTKoM0NRhJyxdi1GTQwt8kS6e68
atDgeCsKpkfEWbg0dJB7BFiWiit1UapwIRhDn+Mb4dkUqxjEnRLHzrfojnVQLw8n6ZTlZlpkzprd
+4AXrjfsNl2xniIeDttH1PC1+JO2j8Xk+c3SkkOsxainQDKofyQcirfgkts5akbNn8Oh4QuVW9+/
/UVTdPKWu/urpGye2/Ndy/Q+ee09ItPe1Vkm+g9jbYv4UZJc84r0qUtLUcSGASUxNRXSiRNMKHqT
o2KAVdi7uvhhBqmKOEigNQongQQFo6R+xFBoTZ0DEd+fUtUH9CvHmBrBcg/kOuZoRBezjE4sK6q2
5HsjHqzqo/ZUe67WnXQjHZTx9T+WRyO2EphGUAYu5Hh8N2K0C8dsP9Rx4lrtprSAmn/4P8XYabhW
YmGt/loedTilEVZadblHnaYlCMu9R6ptLT9qqIpUjwRr0VS2WmRrgpHfJmdGeoYexLLT1lepKeTe
FhQZLWc0NFsgEjNzv4oYSBzh5kvRlIp6O4cosEevgExjLGB37fy3t6m/pJm5fdp9QbnupA62JWgm
ZbferBeH9csybhEXVQyb7dC+x04aj/ZUxOzitXwkB/R+ZAUiBLcHpVN/g1kfkGG5X/zOCyasQJMs
njdkWcX6zoFgnN7rYFU5PQJLA760ZGWZs3bu+AxgbjqlHjWzPmJBzaL1xEILlKN0iidwBXAGVXRk
9pIP5eqWu0ORkfgIetZ+KiIFSkuXyJHOQKJcKdDeNN1AOg4kOObgdDSZIGEzaI44bFsU8KpeduiW
H4nrr/J97gH5q8d+Vzk60CU4t43EE3tX8L55HRwgHraVJVaZ4COmOR8wFIgaRCZpp/GhWsT19vQd
88Kg+PuMh5S+V8jmQTRlsXoNVdfPmlJCEqpRWva9Llrxm5liEvLhh2fYeWngzoDm7kLMvrMbbNXH
J6j6GVSXSb6UHbpMh6uH835cZpvoarBabwZwLgjXFhNK5ovMsMDHUVW8+0CG244lEuqxyO/DFI8T
MXuPucdgDdj+wndZrMeeUXVK5tIVdTgvIy1Wh8xgCVSNJPkIVFNEoMoyMiSYH6+GvDc36L5+PShL
VaK9kXWce+pYZm8td8aWygQKbFg0kIrJKNCNrV8W69/GZZjuMtwhCuM1LM2fgI7wGvaWVcxPSYA7
cgmtX+D1mW3U1cFMn8vjncCC/QJ2546sxzNDt8JchCYcZJF8mJKkz8UQbAtc972s0CXGWxIefKsK
D/wGyjTMzUF+fUwwYqhS98BNKEHhQoRl6VRpKRs1M/AdwOMU8PViKmhoNrO1QfCxpewCHHFOUS41
H2VV6nKf9sqkmq1xf4lBii26xaEbCOV8WDZ1smlUDOkPFT8LhrLHeCMzNm1p/cSAGI7niSYHu8Jf
tKBLOTj16n+VgWOvidoIPtoJ/51sYU/u25lT3IIH0yUp4WE+4Un144CiWMW5v1AnmNDapn5dNMpG
znK8dMcBDuYenbJIvOkB5rbZ5g7mAuMk0SqMDM5kRlhFmZRolaFTAkQ8J8bMsM5YYCUZhAVekvCp
OcRkIp+fWjU0Du+bjbFmmE5a8AqBgqC0awE8kc+WoacsPjYkLMhn/cuUtO848BP7bVKs6DtIF/dJ
Y9etJKvxe9huyA7tb1keaJ9Wc6PtIcrcOCn4jqvxX9WBMYQtu3RnTrj5659A9maCiBKkgqFpi1L3
4b7dwm1a3KHlVyppSdWzqYJccqoaO1PW0hwBxALLydyHI965iLxMppJg2W+Ka87Rr6ny+RhUJqOo
WixB+egUVSgLpWqsq4E14rb31GWw+CQKdBWh8KhjCv871BYCcKdPANilSeUA2P5V2HnWP2tWko2b
tpfeRqFGVE12mSvh+yQ7UNd6S0nY5exvQ8sg/1vKcoFh59Ji8x9wg2+cBpXnStt87YoPSrjJNO+l
rd5nudMqkj21ucDyY/ZRVeCAx0OPNRAYSUzi/KQDJnGzccWrMEDTAOpOj/yjQ6uJJyb5BCWnXVPH
Il2ZMFxw0pdexYT0N5TRxBxYzw41E3nWGGvAtXzjQsTD6eFYVWHJu22H5mEMPVBPuOZ1SbsEzOyp
DC5BlDJlH3l8pBCh54U5+UuAwJQ+27JuSeP81lKvurphY0s4QkFbQ/hxIkqLUYXjiNWZCvskp0vG
KBF8p9a7WWnM4BUoOmtbSF4DcLZqt57zUDXnRV1gdCXosQPNdUASrir8NFBDcCl7AaE+V/YhNdum
Cg+HJhFb0AH26UfR6Zxvacu/GldCmZxFK+UFShlTHhtQBMsZA59fr+xK2NMjButPhOkHw4Z2zSIi
ML02ZTkuDlJ7CtxKS6qVv0go8GdpvY0W+V8wAng/dOMbrew3nNM1FRYlaPXaXoYpcr6qfCcbKHOh
xS1cyIvF6+Nj6y9uTM2dwY9L5cTiPTIcpnaTYmr1Zg45JsACsqjSPbhj/2SQtt5LE0Wohfv6xoSE
AWc5ztTYhp1ifpXQRG/eDfx/TWB+E+W6b7EjQ90uFOw0MMgwrM5/DJvzQa2siFBgGs0y0EYkEuYJ
/ziwb0UtMwvH7/tJ01bTpaxRZ0u6wifq45TJ8Z3SGdbB3lMPD/K4USLI42Wd1P5C5iaEzJSloaBq
EVE2b01guHnqyOhjIJbgykipf7oPnudG0+iarFkw2JnquuFU2M1YVzqCnZI5geQgRVD6ILn25Z6K
Jnlw6CWtNlRSddyuCvnjT3mNKuVOQVHEKoj2RH0kGhcqwRqpcwAWSWrmV2o2cIeKtH8+O2FH6a/u
0+TcDTbjH0L0ycA5INJH0PVf5KbDfFivsAxq2/w8FQ1siUl2IAvYykbMVkiMBNrLkcWr/2T2KgxZ
mttd9cufpkN1hmzf6sYBx+rpxYRstGi3fnLiaeEYikXGKfBVvXg7T21jI3nBIa1KHOQKExKk7KUu
VTS3Swl4McfrPnmWgW8p/s/UR3iroCVWUyJOxuD258Oww+sPbaQUUM0I0yqNo0iQvCg97wKc2XQi
qCWSbuRIEIHx+OYDtXAuuhvEP4Uvb3dViZg4n5mzno/frm7y0wLwR+NyhEjgH2Ro5rYJ7NmpkjZX
OO3TWovZtA8kwfz3RznhMAWkRvpjR/2VBqOj2RDard3wAboXV1N+n3kuAWP6Ao+dpuV2q12toXy3
V5Z2A/KuVtWQcYjkL/gTeEZgIHZHIaV9X1WiF4lCi0DfY7bbci/T8I8Y/AIFoJPjjxSiw/uERX+w
oco4eCwz4GETvZE5e/clMzng0susuVbLP3tTUUulXrHZtNVd1la7inrNEBBe3rNQlF2yTO14z45M
xdo3VySI+fEpTeIpAWB3yv/auAUwVlTUyNg0G5dbIXYTY/1ykw0emphNrsyk7jgMk1Xeg7gUoqG0
rM6CgBBfYxi5znUtQtbNzuYrozua96s40rA89E1X2zkz6fIU1AygdmUMM4pVaH+IwA86Yjk7c0A4
R2gWoZHg2z34YbacSdmkNhYkGZFwX7M+pMUQVXyxAqQ13l2Vpc/mmw0YUqMB7Uqhetx/6060BJIM
KwRGxY8MY279GsOxAoBajejNIzUBZrIz16tvP+vcG63kFxpcV0hTxyn7QsEQ51GDKknk9bTX97G1
LJ2fumlw7qt20iGCiFLElPwVcxnc/bdDwcYKBhKgVByYvtR9XshVz3F34uPS9mps+W5pz+DzCX9A
CALRClBGMshOak5hGFXCOT3mQwrjl6nw3b6rV+IBtBQTRLattNGpyRRGsywhKfg6tyV3eOftFY/x
zmOVxD89lMSoSVxQchT3DYDLODdrwPyoEd1vWy1HWenK32T2Rvw994/bDI2B9fcxoUXWoixNHt74
Njaf8a+SqiuuiMMA8VQqhJBIGI7L7OROl4o9U6BSqgtd07zuwrkDtn3vFqMW3qe5jUKBTfPZgcFU
P+nUpK+ZHmFhSEAHQcbxsPP0Z3B7ZIVd51dwj0Dw4yYbRg5rirkD+O3j6EhYi5X4mDKo91m0Tv4b
L++IZmspVTSXu7k5tnBYSgNB75Y1bpM3ey5jlM+yXCik8+1YHWoN4dZ3mVUfrtiOkAIrvsiaYEYj
PNGJkPbfDRTYKslNuoFiPuGSmTk63jx2QFGSuRMQNfOy6wTitFHCPqqTo/6DCNsjQs7LU8cOwOg7
KU3cpbSZXFAyYf6h87+MYGMzXjswOjMaYgPOLItRqv5AEi+HuaE2YGpYZOQC2usenX0nLd8j/TZh
XiJXyjFfqDNSR0mMWJeaTHCBqYXPiGsGr7/1ZG4X39QNwk9cBgSlM1wYgtOTHH8zaFoMivyxW+zz
6LSqN5A/ViYqCoL0YRE+9cTtpphfmMDeOzR1U4dW9wiSqz9gAOPyv9Eb3DeXlHnDBmzF10vJWZDt
mlOSDyf6Bv3LrkxO1nYBcwgXix4msRG/BQiFDKumH5cLKVdcWTAPC0EZa3PkOLUtpeHP+t9DCsjn
rqnQIqnQcCUi9ueRznDr3y0SpnAkYmEUW5bmO+eJmUep+VQje34SXexnalJDcmNzzF+vHR08bJjY
HmnkJTlhIq4r13gyDiJL39jY+I4o7kVQZg35Nxwe+oOU1nc1jhgxDK9xNMHWJqxv1vtnHoJjDFWp
0tnel7M2hMtnCdDOord+VTOK0rDLll9Ig2yf/FKoQaFBblBq1me1kZV4anbIXBEVJWDfzk8WbQTG
QSQBwgzB9bilVRwApF8R+c2X11yP1y97wiZdfQH8bVhknV370Mq2a+vDTBQXzgrgp00uXZkCQs34
+GVsnvayJaudKxXGmXBxXOq0dRhPBNKmMUhcVkhSbBHwf3SAKdu58plmsGFRYx1Ys0ZSjHpHS23m
d3GKw3dIUU/kna1p4nUqci1AtA1DVIe7Du2l8pkaxmDR+6frVtXFRSqfWPu1frpezrO7LmZzBpEO
nHK6w+YQSJkrQfCuhORx645IzmQf+fV0S1kLAVG137Z1hx9Jq2dadqgbEJ2j4Q7XLzGhb8R+k7H6
710XX87m6aCL4Y53J180iKmXLhB4BOpJ3wA+n4NXKwjL3rgcLWwhsPDfNAWYT1dUtr4xL9rMGohO
cXNjeN35UQNXMK+WF6oX5FllP0eZkh0YRlbp8Kalukw9S9N4IuEAR4vBSRc238c1XeX7wbEi8K8l
5D71d8SlhC37X7kv7O2PYVEiS/1gX9bvr7jYdn2vHhwEOs1NrYSu/hlWARgWwdQb+12yxCuJ4QBq
oN/hoFs57mM3cZfwK7eYkA/tJ166hsEIipw3oPEOrpkTE6Y0EdgwsVpPxI+HrdXlYWeTwnb8m7/4
piBStx6LsIEEy5CZ9uJlJ/rm5J0LBlVvS9A6ZyxV6daEDliLescrbzjm4lA/9AddTM7CY5jGlbEo
ng0dcZGsmsML2f3eQSy+3cQ3
`pragma protect end_protected
