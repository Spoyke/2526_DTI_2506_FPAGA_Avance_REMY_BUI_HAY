`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sqoNZpEVxB2u/j1SYbkfbhJLcrboqHFok4zP53fb75v1PyPi+iCzkaK1h7kn7pEU
EG+XJ22nkaoQVeDbNsh9VIOuM/GDcW6q0Qo0klViOJQm/r41oQ7tlVfo0KVY6of9
x9j8Hk8h0D0xydD7jY958vhAi1uWEc6BUxIPr9gFdDI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4336)
YlSoBPrhigfUP/t/tTuLj+kfsI7cEmqvUCSpnUn121Tug3ekorhewx1jWObgKY/6
G49ZdxEBSWlcOGzvTZ0xm+eL/1iSC4XeNCidFIOv4EqE9V2JNm0GtopjzAVv7J1z
Acwt1AKqEneCAKXWyQhUZZs0SiyS+wAeGoIxWTBQ8kVAZB5SNJfZwl3RA16+vroG
lLpbeItP1JskEplfX+C5B8I0zRsfM4m3X5FdTH7RI7IQzEnRopuwYlWH44/yIfm7
ZXKPIEecEpbsjKRkigx1eZc0TDySUV+a8Mhc5gOF+EXdUH2skSH0rjsPo+LjYMXi
tsoopehX4ARxBoY/tqtmh5ZthmlGJmn6ZGYPHPkIcoAYNDU9XCn/k+w3hPZ8TZlr
Brf9B62Q2AgUq2VV1BEcCAdEOryp577UvTrMAEg293ZVEgoFeSfA8DoxvNzwYGpi
3LD5A7SZM8VRdv7yXH4ji+E/ssqzZJgp8DRJE0g9uKDJ43dKwqNssKp1tJZ3L4tE
R6KYmZX4iKARWpSxhrmRF8V1R3K41amuNKK5BxODIJ74gXMuRFFWCzZwrAw2XrsA
L49e/hJXrfr1p61xvaNZAD7ZJiPxLLpxaIxI5a/MfPqpxd8tEXjlXgOC2yVAFyFb
eu3FtY3AkafqFMG6GzFm658kAlG70yRlQb4xT3361541B8QwP1ski0O1StZIY8I9
kZDWqBBUpx8e84/h8LfQoOlefjeM0fpbxfbiUY9Z8iIDap3eT3iSYPYCEKFSWRxq
JCLqg/HdxVM7ns9/ZDlLwtPy1SzsaNTUJAEIjX+k3YHbpkDwtFjxLHklwJMclu9z
4Ut4l+wpZSdQVgirDjhodUXQr+1TKX0jKbQQ3kCvbJizMg/kA8qNYMF/9hdeACOL
z8Awp3bu9qDTBev8eW8iRFE7CM6OMQ7qzXdrUmkRaK+nfZwgTFsxBIyrIrEw+DCO
/JY3Ln1Ns/Cw3a5HFL4Lx3FJ5+W5u9hTwOXj4i7QHFAQv8zO/7NXWY/9ozNt38ru
tzUIttlF+FwOmLkMp/VItDuAInsNJG8WQMVKc7tJqfPKDsAq+UJe1e9goLr/MipZ
3POnZECrENc7QaDF5K1/mSm37yhW3L2/4FOYoI4VCJze4celgH1aBmjGjcaVDIAa
iGqmv4XTRyDwD8APckHqe40zNg3cbThkhJs56hDtBZdbJnRuoUw2s3WcbsfSM8PF
Mc8+tLYNxyDh6GhoLiHfwPdffhWRzWH3zfxLHw33Vr8r5/vm+gqc/RT8orPaCE94
D8pAKxVkMRtSluS2O9cmTmG7F6p4Nw+Bt5x29bq2wg/6s/MuGWBYCSPYjcWpQMeG
OXX0v6pjKEWZv7HjDA31QDWebFQ/JGQwo5O+4Hs2EJR+KK9+i8IHnHLDD+3beVqs
YgQTz9STbqP4l6yp8mYXq5DeQi3HrQSIuk1lUqRL3XSNp92uFdW+bjT4OYwCQTqa
UXbLGch3O79aq3HCjAO6feu+hO2/IXd8LevdexPDBPur/JjKQQmkrFw6EUPwRwut
zJ4DkYaPx+rbpz0zJUGw1/tQu1LcrNu1ray+xP7D8tPCTKT4fraMVuZVs7XvXa/v
Kc99oXXu3eZQMM+H+l3+xTfRvUerFCk6ZkGvWZg1x6xir+Xqik6/1KbmhsKPw7UU
csNT/IO7EN3uTWL6b2yRcjfVGeS/GDYSSDfo+E2Q+MUnTzHyBaBqOJdfTq85EO0d
uebAO1zC0m5PqYzDOvcL1p4JRXpbwelY5QG3TCAKGxXjmtt5oXzGY8LQsEK43brw
KxVPax74OGXgtgPcatiHmT905ec0o3d44wWeoJ5GKhUkvdM9dBGyoarxxy3bb00R
DcDJksKKkSwX8+WMnnfBoCdVAlweiHgujPU6xqHwP1PX211dZ8jiKjWlN0Je4rK+
xc88L1t8VSIsF2Y6IqZy444BuNqYwMkn1N4kuFGEcE3k+FfafiaWYDBZcHCO/Og0
XE1IX/i6DiPTX/Zs76xhQezJ08TxcgtBRloiWUMBQ7lG4tlj8+6A3cakQwmxz3N9
F23A81kBfIgvycbHsIlO3k76hE/ho/Lzxhr3Ks+lBuuEJcCrKvI+VlqZJ4spevRF
0ptxqGksm83GDbivEQLL/5RIH1seI5yzZiNrBavL/OKBfSoherGdgSUPG2qWbhSG
ECJILdynFqGPXQvXxMhNtSh+Bwsf0JVkr47U9iFY5mQ2bDe+rY3FcYsMj2KHIhv0
8O3glvNsNaEMEhzs+r2l43620D6n6BK2RMq2KfwghUisncuacY6f/B7TTYDI8JZB
VEQP+Ud6AXsVVZ3QHVwnzmPC2s/btXJ/q8/7WDid84hjkEFYJFjh40hBOj+k3rTV
Sodhymqlvg/88vLrX7seqBgV6UrVweowlvDson8ptMXZaVhP1cah2MTvntyuNkpY
Ldew/puzECGv5KbVSujj2Zb/QFuS+OMslSOXKeSDlWQVZmjVRin2zIrRQel2ocOn
25ldwwDz/6WtjdlxZaWOG0Q2TxD3sg/axr2BUMqxpSTWPwqdFu4uL0FsJQRiO1Hz
VuhicFNMsBEAUTxrAGltCEBmC1S1egq58Obk4f60DmFiyXYYh7D7iQk2n+HqxPmQ
ChoN5u/fNikajTohCATuOJFgaNx7G7/O8DkUFCKupbe18Yqy7wprhWgnyP2qagRb
NgkOQXCM7SQUmJUde1Tcy/6nU7jBpD6vJ8o2Tv+LFojYgEhOq+gcFFXlQ4k4DfmY
cYK8gTZw4HwGG3o4k01j8T2PUjIRLGhvnrtpeO44kkUFLhAvQpPQESzE9I3Bx1Xu
2fhAPiBt89xgl3apwdgFFKxIhXd1gQQO6Ibf94C0ushaIATJ02tM59bZye7s4NDz
tUTLEpMU1TS52FrNGUDFxLhA4J3TiBhhiMAV0r8XJWlTus0dYm/I8UISsJ274N6r
CpucO25Hiz7suIsFiMrLeikI86H23FpNPSODgoGQeXtFBe2/tijhDPD3sH39q5En
3sQNE76eamkTfG5Nz3ruf29BQKCBy7mlnfeuvX6P95xISjUAqEBX6a6DQF/9Idr5
AZc50QLchyo+cT4hVvzXAjZBe+MX1tm0n/7xKKdSigCjuwf8irXnBi6glk/kPEMN
0c1Absy7rd3BVs1oRowZEyCi4iB68AM86Jw8Un3LB1VekYzG4RPTZ2Uu3hBzLaCD
IeUjfI8P5qeC7RTdZOPN0ZzNGLbMZVUovcWHgGCKY4GVH1bp2TPTCTAUJZsvuwNh
j14TZxE+Ms5OZzVKcWbohvNBf9nNOHZKaB2nzslEXBDUWHtxwi7MPl0RSaSrKRAi
5uZbIoaU8sEIx+YHLmjgDIBAflUQ+UuGcqDg8Dpdagy4vOPLHmATk0CEK28pzovX
WPS0EuyPF2U7g9n+uSb2BSKu9NZtzbdZuWkt9VBdrNduI+UbQzddR6llkvqJnqDt
77g4P1+UcVezLJw+MIEzPhva8qEDVVMs4vgNjVqo3M76Jrusp1HCjdcZMbJ4+2ut
Sgv+WWPR21ZULkjyFEH4E9lOZM6yLG+eQSOj4VC/QQOw3gM5hPdulAcCmAWGTL9J
6lFBiHpmZJcq9fqT+gRQKOc8YWSdwNIDvNlogtShEnJlBoGTswxmNwVBDsV6rkZY
bojjkoERu6F2yb75t0ahiDWEcoDFKPnw4c1lQShrjqjfRcNarN3EX1BG69CF4Aaf
/1wdwP16idYpZgHYEAJBXNHL+b+olsvbq/G5IxM3exfOD+VDnKpgJsWd+2H0EZnn
Bz3/YZPNuTRg16kdA+krMgFa9FDUDqDs6vC15HtduQj36d0ef0EsjGPVfJrPQOP/
/2f1ehJBlNXMx00FV36VEs/w4bYLTTjErUBePB5cgaSCH3I4ooHRXIziFK8YFhBH
lQpll+9l2qd1Xg2/6zIjQi5DrVRRRvQmOisn/ji4vVoq3IvBJVlypwyZDQv+FO+r
XvhgTFFCwcP++TuwOQAGsQZZo8dIHPFdDsutzIOyn6p5grcRpueVnYRAwHZfQyCz
wak7Si1gS1rgBEd46de1E1oIBiwdHtujgv2xEa0Tx57ma26Vupdd+INYRKOWyK63
hrIdOKZMid0etElPauDXbdQm094JXU1wvOm6grkX0Fw3RBOuja+QPPIpvCI/UJMr
UkLR3FRxRPJQmZ0lc03uUFp2JNQgoXKaKdHMH50+mxvWhI1lOGVJnxhZT/kbjBT4
oU/4afLPPXO/QYx2IDO7fFVaDNqxDgrkKSYev2MT6dn3jFjzcCwcjQaQcC10/U2B
ipopD+DDJQRDZooVV/qH6IfL8qPurdxU2Vn495gitBPdXeQixAx0tD815AIJ6X6+
bYIFSdu+7/+HcwluMvJOEJmdfVbeFJQEguqbawnG03uHnwi+wrKeQLeHlcUEp1ku
JvOPjpgY+WFbLOR4mg1uXJGjy8bjXsGG5u4E4XWFDChx1VrbdJoYN5sXagzgEvtd
Zj1DB6gSAWrbIUr0vd8l54KHKm/gNawVJhKNsX1pQfIN1sDpQG3Q1YmFTsTSG3ar
xq+2k4wEosHoQJNqlSAldK+DwlGG5lIX/NoWbcemMmEEdgtk2kmOvj8Ep7L5pKCw
mCFYOXEheIqzph1XBPJFQCfnsx5fvK8eIenSJEA74rt5acOKrjw4kEVRlx7vUwRA
sHuxs5AwexTy8eyN1WtY0L/JFetwGOZstLU1kZUt3g13mSCJAHG4iu3q+GF9JgQW
YDy06PGd1Erz0xNgIjw0UxcdvLuAT3/L58TrDBz4QpOjVAf2P1S9D56P1V/N38Qa
srMRxGO2NQSeBM+lNjOcoHfYZoEpF1qTJGBJfK/7DuY+FYJ0jwDpqNhKkL50k8IM
OmepdqpIO7SzqUH3Z+nDVa2i/CVyvoWL69UQydTnVjr2pC4Yr/661oLJHU+IkBRr
XRt3lV+lZbyeXm7LSuLoPn3f2zWN+p05U0mH9GJXk2BE10/gbnV9FlD0t4AE+i+2
M+A7V1FPJ3NhVErJmxouWRsYBnbK14LMOrd5SYIoQNkJ2whDFB2MrEkRBPeJngPW
m7mQ3X//BYd5KjY1UHWJ7TcWG9cutluZys4HZqUNs6GKCOA2gjIhTiOWsHcph4OB
APdAtSsRhtFKzzMryXYrfbQX6I0AY3ognr6bzo8KHMPoPcbw9tU/4MFm5hvJaDnX
5BBEUGeeBq/6+Y5oHvaOyXPVU371U6uIVOzsVeyEFHJiEnCJRgf9yUBe+BgOVuZn
SM9XiqHlOpNZfLCafHpWOCwBODtTj3FoyyWTnOHnpz24Dx4LhJBOVc2Q+HpZAvOW
4703KjIx7WbN43dU5gtcnKj2qCK1pnd8K/Q/6aqSkW0vCFedKtfQ278yMNNzUBB0
gaYNe3BasqWcZ8Xv79NinBmB0gM81Ajq6U8YDMxyKtY98RhUGLrP0mx2QV7V0txm
yPx5xpjb9O/tOFVRAZIumjv7IlkiyimKhnR6UWz8k/qn9XB2rD75muBgx00jZ0q/
rI1+P2hD/tHXyQhg2Je06zdI3gh4fs3XSyHVv/wEAgsLS8bWxWCFKILCyFqo1ymB
tkGrdoSNhsX1fDTzyEfjgnWjeu4xFs3w5wM4j+xU9Q0LY1z7m2qd4octYhuPKqgY
qT0CyeeBbCKPEFpo95QW08wBate7ZVAH21FYfLNADiyTuIQD4xBuINsZb6umuYKg
2hwL92O1e+pPls5qDfcJfq2HVA5zxtJYgKB0vPtZla/uJ26xLjA32ubh2dE4PI+d
p8CpGZbw23RWH6ZWY+jeVQ==
`pragma protect end_protected
