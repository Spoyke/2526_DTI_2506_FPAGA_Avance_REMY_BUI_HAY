`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SOWMhT+IUKWLo2n4YvOF9JvQuGdh2mF532IlOUT/kJb0LCPsO86OUf4QGXMw4CbK
WkUQfmKZKUGrwNDIl3b/EFdMnpcFcqoXBS1jPidFzQb2kQZy83YJy8atEwtLztMt
E2CxYd9+Aj4BB1QSq5yQMv7PH44TXGBdCOmXMGMmims=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 53808)
gSf/bqbfCRH6NLJXYEkwS1vTZzxvljLR8qM5Lb9qJ7RNfzQRR1xEoRNkJ2U3efU9
Fd8ZOxwSa1XrH74H+BOtyWL7a7QiIwQTFSX2LDrPfppkrIDjpYFE6iiyQTms/akz
YbaAfmw1T6xPwGgpuCQuUAWnHomtlWgUSdnk8GMfL2IzzKndzzznfhGy0h2Vkizo
ZFOSbaZBjPVZK/IYohu8+/jUKgUEYXoa4RyMkeG92/sal56ghwrvmNAJynSQyEg1
A20B3VuJk9Ed2GQPoe/EhrSd+GUOXc4h4NcAl/Q3oV0F/z+7EHyoC5W2vgkM9nLH
752uQ0ft6WIh5rGQoN9bUWTGthavSoSpKMAO1Sn51hQmepSyvxjlZoiMtbaN+ZGf
a/bdB4bPeserDjP76gIE6exMFcyrfWZJYfmlG6LGENC7yDmaBeA0EhwP6OspfMn0
iL++NvZ7kKIIWynM0LIrksttz6c9K+TzZWtld/1mHsQ5C8r3qRwQFR4V2FlZUplr
qs7wvONj16JcGt2kHqHg3Jot9USCnvRE/hZzLy0x8krr7fMy4jF/ymSOIsgjcxvu
Y6VHr9nbY33eaLGsyyeCmdqqVpaLcOpgS4WRVBiuIr8v/ky4hjK9SbMdVbHl7QIv
4PDyhURakRmMnsN3E86ycLO6rXGT/Yt4Ijay9O1Goka6FtN9K33TaMk9aFHEN5q4
vOpBHsXr5tpCt/yp6YZ9d7ae9qyAZXkICgBWKtpaVaLBU3YiovnPGT9y/+7jy2AD
TsQiAwl/SFMRjUKSAx2MlUstmxrLYuOlTP9pOrKBcDmrOz6IeB5eV1Q2U6gJfyE4
LTy48OCiEvZh9U6RcecYfCYdWpxkc8V+rUBvf5bTz6yr7H+BLvkOtL9YRwj2Ggo6
Ed3TqujKAehKa/59R8PLFNq4KTxqZb8P66SsM3/0jPaBV6tR9QGOEAWJR6Wki5OT
2Hpyb6kZCP2RnBH1esrq249wYesM/CDdZKjrTdHKtgxgXtZ29gt7xEPiNOuEjjKY
74raWJSu5TeTglgciMin7rxILMNVd/6bamiA06lJSwN3EANubL3m+uhXf63DY6h0
B6MHKut2K5f20wd6eQqT01Y3Y6+oWVb8eLbNUU8obEhKPAZian9IuKiY0W5kdmbM
dr3DK+FAnIz88maLwPdOy9+6Oq46iCHRfqufFL9yZ6cE+st4GY4wyM6uqhaydOIA
LhdzGURgeP2gJNBFxxqklYqe0hU2AWp5ZyDPVTiY0pS4+6h/fCFObrHbBNW934u1
q25yuu/bQ7bsYV7WkOcNFiR9aOiG+DbXDFFAAnYYJs1kKZS9rX7kGXYPO99qwEwL
XrWBC03jYyzkCUYL9KVN07N9PGLABEFZN91QS/s5PGeNWXfA/4wR8fo3bI729gwT
wAOc+Cp1EVKK3yteDuRZ6QoQnUeWK5OqWQQf+mHMiwUT++OR0YxSWVLae8u6SHvU
H5EL5wQowtDf/rtbc7HQiLb6U6NflAdI2ecPywmUuC0pjbwpMh1JjXkNLe4MC6In
6FfaGM9z51weaeXPWgZUM+nK9/dir8n7/ppYJWBPkqKnSyAKShDIsVDOMCTjfRl9
sB7fSHo3/GTJCXbmCkuGy04krtk8lWtUm7bkmorvN51r9Z7QDRPHMk9++jpIVRAm
ac08LaqHhDh2vXXwRUmmTp0gxJsB0sxNkxRx/QYraWK1dPGtw06HdyxhvRISXrdZ
NIrdDh3bmd7ta+6fNmI+IGQaJYbQmWwNRi5F0sC6ALVdeKFxSuifhrjVza5Ioltq
TPFSDjLl8cyiwGs6kABNFeMFg3QcV2xEN+HpjHV4q6ndLMd8WVoeLzDJNdYCNep2
FtPiuuiMYrCWKIf2UXOci/g90Eps9o2JPj+logyVzI1NsixtiPmLpKELRJXOm671
QRf1ywhxmNcCkzqTnkn3W+aNvl3Bvh7cq4wjKWW1250+ZxlcsCA6Z7QMZwMdNgEQ
VQiOLrIGBGaZDcnG3zKDUU6NXadRHdIThLA3T8wF0g16MP8y6vZ6rWCWREOU1DKT
JtrJyhxjI7ynCZfJ4kpivCNYT8BFXGVA6TC/rCvZtCUHCJsn2WHGQGZFF9Ws1zed
ke9Z81pz3n9cva+/p/BVaMAunKU7rnz8DTC9LCa+kwGQXWllSX5WZvH1yt9rrJSE
q6gxED9RA3OsOOHDmtQa+UXnvsLcx5+5YMxRdOXEmjcBLq/cAIapLPuRcYmBPBuN
1diiCuf/2bpZ7LqZJfXNha8uwRAM6ygoLSLryJMCXo9JKIqAbT0H/6D7pSLplZla
EzU13frirtP2xcLgD0itJL3IrB+bbxjPb4XYID4YNaCDIBuH2Xw+y+v2c6sBhQVN
FHlFYm/+WDE5P0odR3ptcM/VYrbDbZJ6Go8VR+bSDGl3PB1tqW0nj7MHmhjILaAi
favFuoegFoVfZQprJvi+WstkbedtcTWJybk3495hObJeFCJh1KTmUIg5P7QHKiz1
xppyTEI3CitWjY8mM2unJ/4oe2LbDm+boJ7odbFD4OLatX0c3L9V2zeiH2be2+TK
ic+dBetPlRL2v83gHt6F6Npm26Z3fOQSBp3GNHHy8JhUpZLcwNOXNatAkUyzY059
IvQop5o8k0cRCHBjbJd+CjzaxY9EBua+Yd7neDbIWEjcKdVhE1vY+VqdnxxDML4I
SapWCsLn0+v63rgv2UuwSp2cthSWicscwDxfseh3FoKyfKR0RDNUiC3NVUf9/uPW
h40/eK1SCBM2+tXlXGgAMbG13YkMDRiJBt48uvo5fC83+mXZMkKPzZtKtUkNDUhF
QK5mSAb8QILx8RMkVmt+OwT4s3huZHNNeh0vE+UEz/1xjNZqWseNunqdFuN7evQL
q/OEJ6ilfiwZdmekpbThtBi/dak+LiBG8hvU4HIoeSzYd3S5mVPNh8aq8tnaUSCG
4eW9oIraDTbhaD95B9UkbqEgu6E2vWyKo0GguekbXETteqcRivI2QOLda3EmMqIT
+t86Q1AcsGTFv//yIcACOJIPadZD5PpW5u5BguVYyK8fy5jlw0HcLSWl8nSqX6fp
NurQJdHtR36UsN5YK2MGngpuBLb8L68QA3UciObIMMMoGavuzpLY/HLkJwMmS3+c
87KBAGmWe87t1EyKD3ztnjw0lsN+nrNiv0pBNrcTRXuXlrC6X3FSsJpQuV0rODTR
EzLf9+/Drps1njLp9oJkeiTG5uat/TRPUmAdFS+sKCRXAA792HKlt33K8GW6Q+QY
9/FDGCKzVbUFpPRR7nX1W56uWCc41/Vcn/L8Kbn9nOkdH7ITPQyyZSqLkAY5cEgj
PvaQRW9340p7tCR48+LW9vpdg1IS05y46kylP7/xwAVfD5f2MiETM+A0XZrdiveS
r/sd5lZX4H7z7s83giZjwGoER7XS5ii1U3Jpd3bT5cOy7oSKzxOCoWBOynOP1NJT
PfeCSen/LiuZTInfoiHIGDkteAp/lGx2EoWFcUPpffEzitOOZnzlfWcHKA7YZ1+/
Cnmu7ffdhv5tPWv8cTL116/5KVjxorhzuWzaOgE0pRioWGY3cH2w4gGqmc4GJwbt
HzAnpK1Wsd9SfYLwhKDsJMQ8KwWFv3F0go1x3Ci5PrVJTNKswrSTPkuQ6h2JgG46
oDdgfbcyY9gZlU/qXFSXjDb3RP80EnTE3FjEgCnl932IDDPor5RPocDeBx0bS6YI
r2Ctmw5tMBoZtui5GNxqyYhKmBGADnczt+jKzsbLzADE6jY6T4o+h3ep8HNNjpg/
3u/0q2I2x4JryNfZqjzWnSV/HzFjRk1FhVADLlWcAopnip5TynEAS7enagPgUhar
UnG2MrwJrKG+J6TMyAquejuHivaVj2yhCMFreOWRiNvQxZRJq9NI+IAdQJpkbdcL
+H7zlsjteJiAYESIpdzIAldPpoSm/pSUo6PEuKI/rIkki3q42vx+lmLVM/j9ywUE
trlDfRR5WDB4jOykiCHF0CDg+bgmPcrGbPaBHSjkv5v/ZWkJzXs1Vyq5m/l60/Ei
9e2vh5EiPpMLnfs9Zunn35VObkbNQt/ds7gKQnAPWEBClp9oOVgaJ40MqXaqE9pq
o1We3zW38F1ZWHHEdk8LNnlurZAbDAGG9Nc868c7G08Uv6grn6iQQJzU+TdDlS5h
fxKY6o2pQ+ZV3JJP9x2Yr6+s7YqtAslgJrglnHx+KrDiOWYPO6DRVLUwmZI5NDYm
QS0fr/Btqo0WGviPvnXcqSB0LzoUqutbDXdR6w43j4ZPqZHKEt2rnjoZIX3YRh8g
yUu3dZPB/ka+FhzRdZhkc+n8TLYPM8fpmKtM82OQeX6WVB0L0cwk3O1sS+QY4/Zq
I2K9/plQ73nYtHR4Vid/rcJv0j1INxG0MJtoJTHQQpKEdBYvAN2LskH5nsSxPS7N
igvcO6oEeEwgFHx7gOBzPAsiVo3AXGfwFJE45GvvrouymHz2Kl10bKBGEc3eYJD+
1C/g8mPtatb5m0Nnpf0xRSZzY0t+GkKUTs/YJs02fe1FGWH82M2++UfBaaGZPsC0
HkeUgFMN13nn3L+QgAt3EkBVdVZ2WdJpRmyV1un3B2ed8DspwusWFpX8Gd+e+zF0
ZLnAGFBDZjypYmkhB3RypButzyq2kuijm/CXTYowWiUmOLNDf4ZFcR5p5/0AzGUK
ZQ5gJ2SvH7eRkD2+8dyrbHcHdcx9m6HgXPsE27pGSW/EcPLypbfSuvo0Axy3VCoc
M2FdauvqOW8xEK3YCLJNUI5o2cVMmSiTxGzs8k1BoEb8Q/ohgQRopjIfr8zi+JR8
MLv1t/gf66JqwxA69pfXtESM3Ei6i61ntfR5AxNV47XTWnxILVth8YW0J6RxjuDz
jlv4wiM4aMNBQlzGTFd5g1rWpVJaYkrc6JseFj2rxCuT8Np6LlxuvcGlQs4/Zqu4
7j2nYUYnSBoutzF5h1htkE57G8wmcbOBPevrcQIjosg8nDq23f4TSAWiGOd0Px2s
0G2IfFmBrJwGpgbq39R0xoELltgaN7wcrBtw8GA31AXfZ7Qz+CEmtauqMNhADPA0
9AFhIXsVQMAYI7HeIe80lLvbansBXYJ17H+xhMktMNMz5Zbu2zQs/CjxyQ93tZlc
0LautfgMFezoAsC5aCatX/R+f7PGHLylMUV82MaeVG6J899a8OR6KwBTE324epYY
pWMqKxIL86Pw4D8JqAKMDQOtg9H2Dr2j7MIUf9c0QSU7v/kRO7zlmFk9K8R+tS3K
S972lXKrmIEJR50ZhJGwT8S40LbDDfO91sYU4GVE9aIKNgkPlpcVNQBN8qeNIs5k
fJr0VbY7AunkmIRiM/GwYv1H/kJUZPzESM6tX2TloBwtFt2cr8Q25zFkdBWDiF5b
QEXCTu7+glhzpQQFwdRKdvDtjeSUzjTQXI4zsBETdlyOeXDYUnVXZNCrequLnK6w
G0yrKHJZDUDqcVRLcqpauJnhflmdvsaW4kxIZeo0LNzgwfqgT2RSBnnnARsAR7yB
//sG03HRLvwMWXswozPn5Ym3DFzkXnZRx0yLWybJ9SEH11/tV9UVY98CioxIcASS
lSgalE+bOPqqZK3PX47lCuJ5ezn6ZAIwcbIxxsqVQRwW2yqd33x6zPmeczVHKMLC
JnvDswsaWaPJAjWRN10p0p3bXUmmt/4y3+2L3vIisRN6SSH8ui1mLgof0tmKZTMM
bR/78IEGWRQ3REGNRsonAIj17UX91dn/DkB9iA0w2UejQq7Koseuj9bLua9pEj4m
XoCjM3+iOL8+aURUB8A2gPn797aaNzmaJa8B0jdpm6SNJhj2VYSLCoRy40kcoLz3
fUQzKmR4E1If8ML/fqZbxY9WVPq6PO3A9fgp0ILpdthnuXArRPCmgrCPbehG40oR
SZyP6kbcM1MJQ7qbrgtuILMdtwEIbdb9j0G2q5WtoVGwl1ef6fjpos2R1dlzQboz
LyeKdF8+s8gEgcPo76xDAGTIDZDY7M3h+T3sk5h7RrBJD3pTadPCdpcFDHGyszYQ
M81WpbRwbC0ugMi4tk8S6NIEasrnGrSNqvkpnYsWV/Mm34VlYXL8b/RaOh1RXDIQ
xgBHY/crIfgnVjAqAMwx2jrbmH5Be4862fTvSfaJQLeF10ugT+e6Hn0M3gbC4vTO
dzA/plFoXpxUUHfaLvv3ri59WkBNKkF5XmYFmAVqlytDSqT8SbUAfb9bD7lLmRdO
+l02ikd3g92jfzLZlW+wAtgqHwfd/M48xDeeHCE7cQMgaV/AuLLhIbyEUqdDTOOG
vJgOICQd2ptPoTq7xjJcFc16sz6uSDnktK6GP9gedYXHyhwe/vMyjW+HxGb2c8GU
6sIt0H4QHooaFw8H8n4TWT26XRRQJHCKAwptY00dpQT3osxNdJMl+5auOeurNIo+
F9xMTJgo4FindND9oQ9gr6Ovxm5fz1a/drONNHh+e/oT/YgEx8KMW7r5tbhT/BgZ
F6gLlCEm6CsyHuHR5BpeK9LwzVYieACGcXYHsRS6k7nN3RCcjsy9Hq7t7CekpB91
+EtGcTG9aDZUpxugvnoAY+rVHX6XaUmBGYmxnRFLtyLdyV9E04esu8JiIGE9VMzR
pIy9gZ2MVCgPFtN1uQ/m57cWxWkrZfbModYn1Te5/WH8OixVSE4T1Me5Hln1gia6
JIqu4AA7TiXJpR309F9M311w6wBP11qPgWwfCAmNOztuJOvJ4TQv+d1Qj8joKqT9
VF+rYOlltm0HBkJJ8aDHRL0EDiN1rJf7JpMQUvVX2e21rXG8J9FJZdElSk6oSwGo
5dE5ur2JTlz3lok+HYkHM4E5FbAZbUG4g15ht+XV19mH0PaJus9sxc6Wb8XDyqqs
1a325Z8t09jpgeNmNOK9HRc98djHjgw3Wgd8OuOU5DJPnl65Nix60vZcPnhnD3mb
agj5W+0QszJrMzB/Z9Ex0v4iW4NtcfKoQ0Qix3X5zbf/xQLUtH2Bn0PYWIrzn3NB
eMVjzsY/yCSFWnqLjIJ0bJjaVz+CaUSJOuBbY7f4XOvHFABCVR8UrTbMQAh7jdSy
U0riYvciTLTNivgWp7VYR7M1v87vkIM+TKJncOCAEdT/VZYM7z0tNjbMxNJCxom/
Dv29pFh/9vsxl/EpqmxxXjgKwgWy3gbmzpwGkhqblek15f3bxK/JmUt2Whsus13b
t7pdBaBe09npvvg9FP36+LWDn/STUn2FMnoQrQy+tMSwdn6CzSH9xXiRNUsFwUnj
jr5ZKf9bn8ljaUqsk/iJf06Whr9cEgrxm28SrvCtRz6GQ2cVAt23kTagg/REOvoD
aQpHTlsFTU1L4hr2VHm1vn1fgaXCgMaBXGfXAom29xoYzS/9uH3wgTW1hqvGStQC
BA0a0I81lrmvCQYltZ74tM6gmbYsABpr0okHrHe+1f4KmgjZ6V2J1doIZY7mCABD
7NOCKLV7muvdY3Y41HpQ/WHNbz8cnmn/SNTqRhdu+LVt3fNcdHx9TydLV5hAGq1q
QhuDtDhbmWXOYQgDspG1ylZVi+l/bUTuEnixLjmBsn58hSb+9WnH2xZwRbllkcTJ
+PBWTcQ4wkWLndCfmTqGYnCuzbBClq46Uv76C0aF8kX0n5TO4uB6vJpcvozhWfcu
77noXt+5YmbNXWB1Qm/omT0EKw9nM7at7YXzAeAIe8BsE0n2y/J/EhGR2V0aEAY5
rrxpzwxBfH/aN83MAV0zRYNPSFHXQOwR6xEmsxq5/I0NPtN7E7WtwrGustx9oKgj
hsgcg5DY7P42WZTW30ssVHjpRcWxzToE0MK6xPAFNeJKmFWp+OxBk04csGv/KVqz
hgSASQn8sZjjn/gE5TzG3SMffZR0ztSLXxIaPZ3mZESS72BbufWivwe68oiSL8HA
t4aBThAsLZPabTWlsA4X3rlEF2JDfVi9L/5qtADNnI9k2vV3i5X2n4J9zl3muWUb
5dKOgPCSDfn7uOI2ULxsWwBrCR43ZIuLmfemVpQeyzVFTqsmFjkdn0GOaj7I3Sp4
jPDVZ1Tvw0rfzSpWtAm9plK5evHOdvlNkxFKFhu173ruoHrVR2lGhvXaZdeG45ra
7Bu7UqIyY8WCMBOXONgZsGOCDqe01IzEDSN6FEDILye6HbBMD0s9rcchd3zfg3rM
7QQ2G6tOvqRhqT7J+o6Y1ebsY3YbHfx5jwUvoLUwBa+YB9I9SsInL2rpVYP+cmQQ
xuuse4ePX7W5MU1ptUEUkAeBOIF+LA9IW0OfS62J+xfgAvxZVSIFicL7q7aDfMLK
BwkYjpCyhkchME/3KGrwA6+cExyb2SCb0/hXnO1Kv6UPYldmGLI/Z1b2Xz8GvQMA
ERrMKbENden51Ya9y3unh0K74NVK/BvLPkBU0tXZk3BxRtzRDZLv2uShJRLW64lH
Txy34KqFry10qhEaBf4mVLJzpQzV4chaxIeLoxpz/+xluqH0yYDNtQXoX7H2Asze
DohH1Pts6D/lfsPWb4QpX9MNcTLLGD9vi9KUZEmgZzTXk/Htm12vRwfJ23NzU/m6
btrGc8wVqI5irfLtcarw0Z8bYKmzElEJPBn6zlA5WYaGKObuGcK8oCyycyH4wQx+
IhTEzcmdPsmmH4EAzvJCuxK4c2qYWSwykin2xBw0KOnPJ+/QtKwnVNXsI4C0wJ3n
FkD14jMb3TmjU0Fzit+2OK3jOEc9tKzKHqiF0cTsW3OiZRuXqe2pqpgxKId0QsCV
Mytlik426+Do4/rDCC/NpIVWmaQsbbyMTW3QavZGrkLtKc+Qgoerk3fIykmzpB85
tB6GWSKNTOUhiojExqXRJAvVWU9N+jFmnFDqaDjMiKt7wTjE95C8YQz+LSIYcmgc
sTT/ectEiy8wF5fIxEp8SQhHJRyFVKlGgqduM0UA58C7lEP7CcENnqAKrRHoKI+/
GJ9GAV8ewtteXgsn18/cYprWkpa+lF5pmVW1Ceufil4Yo4oGqA7wVUDjdWpmNsjn
DV3K11AUqC4PKe92sehSsZA2tA4p50yiVttBfhD+Q1QTVc/Sf1xALYfisIo30gxx
I/hzJ0Rsl5Xku6soq5DntuQRqhe/lIp7RXyWRisKVVmia8JcBYAj8iUSwsyMhkBx
qD4VxcDsskUOkQWXK7LIdcrbYmc819/sYV8T8yAqvciknlO763GPE17fbrZccj9L
trELvquwB17CNRLvmj+o10do5k5YbTHfIHGJa97fwGp00bmrcco6fvBwfaXLyJu+
MPsduo1/dfgGoqPocN7jIP2Zs2htG771Yx94x+w0kjLDSJ8qHguKB0vNDFXBchVG
q/K9C1VP2O64zMtqFtuRBXm4fP20pzweQOxmYCci8CTjMSYU/NgD3Q65RPcRmhFg
R/M+pFgF9yX0YJ7LL9BybHyumT4uI3gMwNmk3NthZZifS1FlFzaxX0G9bfoN0ZJ9
OPF3WcAVvRHfkEo9QjVaPSx/ZoZdqMB0zicRU0LTyPIR+lz1sZfL8HJp8C5PSQ8R
Ve899gmhWpL1YhneUs/O5jruT+B1HmNys5+vrM8tqxoaY+3NIOhDlZnlI5ZP7qk+
o+63ax88cb0iyODpgy0bAb2emttZMS5fc7eEsIoIpXYYnt5KzEeihw9vRboDHJjG
wDufE6bdgye/YAEB18kfxZYZx6I/Z3zuLGqXWqbAaGvkY1Rt/vR/zNBwLg1Mc+Y2
QlpMFhwgEL4C+lUH+4TCMOOFyKQoYIEj8YfE5ApIWGlckthsvAUnxDdS5tKX53vS
vYqum4EKoJgUU/AoRqlj0yITY6U9CQOLo7SomueZ/A3YzBXJ/gR0Wtfiv6Zn/VYo
BqUCs5WgeUArAZlXkihIs8jyyR1tx1L0M826pwshKk2KarcvVYoHJDJ6uFgklXgg
XqSZBDuVF9xmd7PwWMmCLICuTr/ucNj2hFSsbmLkdUDRso0zly648qZDGEZDNiaP
f9OL0ossX+RhAgIxdk7yobb0PthpRMackvLkP6m7OyETiK8KlwBUQ8sT3SkqKm1v
Wy189bUyhI3k5OqsQZcsuVJR+n1FaQoD4ASNoFf81fkX/InFpMNOKHbY+4VPXQQ8
F2Oao5Dhts4GekCx9pYS3LD5PxfqoTIhC8u9swEx4qFq1D+JaNQYN1Q58ygN4ixN
gY9ngCNAFWUqetRANVexTYkJD8htruVFyk0SnopjEmigcq4pbuG0ZvDCRmD0ll8E
OPitTfYPYMuDIituMJPycPQT4Aoy3oi13Bdy6mVFOu3pm8opIQs/1UTT/GF40/Mj
0grsF+Pgwbci7Eg+DZcr9hof7WPXhbZdUvW8A4yXpT0eEkZW41UY71k1Lr3kIcCm
vB1PfTSh7oRptx8Xzm+w35JSzL1dUUz1/2fjz5iOMDLrDUBP42+M7zVUe6o8D+d5
+i7jjtIYZ0JvbTGji/kHrUrRG3qlibr8IK7Eh3qXR6czkptvS/FjfJMHWNtCmLko
Ayi1eovE0m2OoyHlvxrEpGjhiASvl47cYXRIicrqnrlHqfUQytXaT2dLOe8/IoIr
taaXP+lRI2eiiad25g/57hWWZWt6Y951UTrcQ3BxmrZbuporFyeawwGTYSFU7t2c
iX2FI8ovTb2MeH+MYSDtXcynYgXUpYnm3KfUsPeu9FFB9CDrK2SqzCqYvuGDXouL
1FqFjSvdnPkWrbu0cxqJaCKcHB9avzhH97Zj6OANseHpAkGYRh/LvmjyhpnDSfMR
+kN+jyGm7a1ADopeOKdcX1oegzYRKmz+vrH5sdEPxAL8pTFAJyWg5UZOqVZpT6LO
8h1HK16Gyv422IQRHZBMJuwZG5ueDYGa1Lso9lld/iHUsWb7ACfmVRn/PTI8W57W
cFVHWgWzU7AuheMk1fGN8clQ73Oh2culbnaIKfdDzoZqyZtS91CK//ZC3vBjUPB5
MUfyED04QB7/e4mfh7OY4Zbztp3ViqtalsVtZpTzhyNHmWBXPskgRjVOcCpnoK0W
DOUQKssQbFAUiPBC7d8jwjtWayHyIMzRvlLZ4Vk48sxbOpv2GuN9JhRCiavws9i8
2fSbDPz/cqGxqih/F1tK0XgC725/V0g2VQrJTTaqyqQliilRN3ALz/HIxVOZai85
ghIQ2dYyWKkfvyiJCLO1FINhxvOUeW1gOoKtQaXG4eIzQuSaP7583T9YtAp0QJ4n
6crLvfPKUp2MMycc3BlCm3ZuewB4BF4225C2yTE4RpJpMnPYOFLi1pshDeTEy19m
r31b26IW4xMl1fmSy3vJNA/Ev7MTbBxZrtRcX0CMFV40M/OHXUAv+GWwLoUrdYWc
3H/18KyyCR/z3kD74fqfxM8/oA70pU1/BUD9ymaYt2XrldLclDNhBO6AQW/dF1qf
Ya6+DipTDNot5ORgF7VRlwH7buFcjhxMA+ab9LFTwLK95zF3ItGlDIeGFmMW8Hxp
jOPWaX3C0z/3LlGwFq77AexTGt/VvRyxLI5iXnRL/OE/Mql2S/0C3Zlnn1BfEHFY
k21am3vgwo/3h5MQK2jYksXzWAeTT0H4QJw9wioOAkyakcHu5xwxvZ9xXoIQ6Kdr
IfJMxCdf9rkBuWOvj/y93CRdtTwmMlwroaW1M+ECtoOlUr6BqvxGzCB+odpRZ+wc
B+qet08xuaRwmCEZ4Mm3iQHqjL7BRNOpMrKQw0DKmfuN51p/umEUocwDPjVUEGcJ
zulyGCtFLv5ii0r3T9SttxxyQAeEZ166g2TNbMW3YkfLs1YzB+Gej4AujNP1Oe8C
rwCJdigaJp3pMN1WZ49tBvmQiOjfM7iPoWDrS6+TaDHUW+UmN4UAR5AMB15UyF6S
S4vuue0jC3ppNRZrwXDf3Ye64RAd22fL1m26DMgDza6BCZQPeBUUEd14uDuN5OaI
UEX2wl/gpzlbcfkwCIsQFMRpZxx8SwTPTGPgTZ6OhNyLtCCLHUbbYuy4CGNDo6Is
9i+7KS5WZ36JlOGnSxiRSj2eDUc2ejJIB/RCn7muIsN6uY61WBVVN+WJljmKUSYn
NHXWIHBqYYbBSCHt+9AEdhytqssLQ+rkW7lMtEAGzj2GdoPsdOyFlHu9rDcUKVP0
c+tqsu7vaCkhYaMwZW7rIfW8FU0C/cyBynI+dOB9L19s93Cyhq2BzaNE488Rz+vY
zrLENh1R4c/4ihcUj4WyV4wcHipeXL1ggNHfNvM5FPqSG2/EKWyt2A9V6xZClCOz
WlN1tZZRySnS17a59YYMyTKtJcV1Aby9vVGmVBUxhbBw1Rs0l/Uv+uTGe4OrrY+X
ytinNXoA13WlXqmP/f78M8B/gvQ7vVB1sCvfPaxwnamchiuG5OUTxDxApB4DF7Bz
9KfgvO/1+dqQk3u3aehGIacEnW+Cfzw6ZFcFKQMYH0wMGaRjc7A9807zcFUIGyYG
ss8tLRTeQluH95GraPKfCDL/zmbjEohiGADSncPWX2pPcKKanSka6hroq8/I6xmq
3AVeC2ftR7OA+WLDDnKzdY4kdkRoU8mXOtYPCjVLnuf5ipku8P6+ERGYLeGKAOwQ
t2KhXsBO/qIo+ILdO+EbCDF+RPDYmQvOjbrrK+uBNMZ8rlDvgE5M+P3CqFAeCeIN
tjLjOsshpz7xNoLIKqTh8ijCZUznEk1VdxfKpJg/Vp3M+hsUjxDaJBe2IxuBpHRh
GKwkre02trsmqAwjZ2zHm2AspWgiKcOW4UQEPltf/0C6St35jmKLSwnwC/HdPlMu
9+9jXVhNso+YVja6oBkHAfS52eUXQsitkT+MVgkuKIKLLX2RuMfRgYrtm6BZ+Rkn
Fr+WZc8ULS2vfaA4h00FV+Z29vlc/Vi/rV+vgOc99VviZlNmuslCW59/viw/VFoh
UZo1NtP4QDycdLghTQ6AONCDCS957NngD8OTyaaEVGRm2EbOgnHuLf6rMSWR8ZP8
jVV/UAIHZmAjwZiqNx5pyu3lXSbkB6YL7vmg05uTHDBJkQhcradhNvwXUGH5neNg
zUxaBPbIhVOGaqDh1CNUlmqUE8h027UTWJBqGiLGBmHrKiDoGfHAjE81szKaLVTh
n6KULM8on6R2K06VG3+gK+7XlvZIDxJ2EV3+md4HcFvY9oqj1TIZbuqNNi0nr0cg
KlKhpVWE0RqYlzISTQz2xEd8AHYbdK/+UmpysYdWz1nzjk1XfyEWGbR/toMb7sVc
sdcBAdoREe8XIXgnZ3044bWVTAxEA+0tlRvYzLgwxUMyeo5O2FA9HxP2ThN3mFc6
j0Lus9zIWtRK+NtPJgERuom90l1EPSoOn6/ssDolqeBnPuuCVG2M5GYQ7mownYTS
TRllRl8+RDOSLeFhIS7Akg21HWLC9FvaN1ABpdbh70AzeETSgryE8e/7sHfRVe0n
WxhhhCwLQJhuOLYMyBvK+W5ZKF0DgpxMnKJvFkQRt5Eca2HAem7ht21WYhqgrSar
3oC0cx+SqJuyaG/cdESVwmFfBO8ECn6o3HII7AYJnxWr3mqR0QG9MZr/e7Tn1kg3
gDiHT/HT2v5tsoV+RMTsoteHPwgFyOwPEySQzab2V1c1MZLFwAEefNMD/a9FpUa5
nyRdrl3Bl14D95uGNau+b+ByggOKx1uNPeTcq0l7NQw/DTGGY91GPexR9El9B8b1
Q7XGewXw9BUMSS2dPFmVzqzbr6qmm5Fvv6KUk6EEGLcxEOhlHvsJHIXAZyWGWO4B
APsZaPZlOKGbM308TcPny/yFxKKp5lcIkYOehiK0gxJ/UcjzIMQllPO4deiMwovx
9XOAhS5BcpCAuN90q3ml/uyLA/+//KVdlXCCZV1HYvALh1Xm0wD1Z+1TfTKLDhgl
OjvYoMWaKug7103AmXiFiw2wWFrDS+UV/md5qF15OKWGbSCsC3SLSqmNrxScujx5
hmRqqOShQHPPkqjJ2mncKBr8tE4rkTiYbIizcv0cM3NYjIe4p05OaBvQYVkL+clE
njpPJEzUTH6SVDZpH8PVk7I6uY39JeDdPhwjo/QxclplXIoCG3FvbojpqGIyi6Ag
bcqW7jphwD5kVfgnQHHUD+SWUz9pi/BCeORHlI/ktDNzlWYgJ+HIg8y+uo7ory19
/20jCwrhKS8RrRVPOxxHD0ESL954oOSCTlAkgH8n12AgarxGTUNUlrk+6FP72NuZ
H+ywruuzLqwXbWmqJrzZob9GX0t7wFaJYFC/y/Mtvwh1xzzSkoCSHQ0Cm7IVOB83
GUjiQuluEmLJbJ1Plckm8My3xwyZLaUfsTVrMWOy2x3o+IygpAeS/nFZogkR//JF
xaicEj4XuduVsFWYzWNypKV6ABzmU5GhsUUQl4qdE0vRHUBwGYGZBwvvBI8exYN6
mYlT/wmEPdn+ymJ7GXWmv2H1AFUwBDgjhqW1kh9Qg68G4S830u7cfU8mTOiSkxtS
1j4RB8+DZXjR4hOMBPwbtk7r0Q9w34jlpKXIimf6eaTOpeMssmbIYvUT7ZPNH2db
lbMEiLetGAmMR1BUcwIQcVv6adVix+ywiP3JXCN5SQ++wPf5r03bNRBfn2KS+CgE
NTze054I5o6U4U5zTHJJ++xoDGRanI/zDKGDReWy4PX9D8zkUAEcRKFZhXpJdkL5
faHSrAlnFueGw1Ng7NchP7mtPJ+k1mBbeKuuF7dUu9lrdy2OGuFDRvSuhrHFhk1X
rqn/EOkdcLdCp9RgzmZ6cTxOf1oz/4qB9J/KX+orJqluBsHuE5r8eV+1cgq0LYEy
DXS1a2AklHn7O7ucvI4jnQt/CJWM4DcqgALYFh11L2i60TBZ4KNSDu/EuD6xGc1z
CkEdEGGFMBHzIIp/WcOntUSjwKTzkOAsGXfXapjFIM/f0TvXj4GklOf2Np+KAH8k
W0IYMGbmmgj2F3U/GNqUXQx8N1GaDnvCvxnhzybh22S5mcuDyjuwz6xNfd5PKqgt
XY43hyXhyFOUha/b4guy1GtVh1WHVxKvhzWvUfuDYjq4FHvPFxTtk+JvKc2cwjTO
W+ve5DywavG01gMHuHRGQUGgMaV9w6dVqKeRfSrYS4z3erR+5DHSN+byzKyEysuu
x5eu+/gzQuMd0Jq6SRpPyfFQthvv9c2UggkPhaqvuDtKCyR0QArPNeeE9P7PLemo
OG8B3KT3mP1vmMrPA9X4i4X9iVKm964Qzvllly7mdZ8tMbcpUgicYdMi3DwFpcx5
rMk56yJYzxKeGxVdWD3ZRASgGH/sX6P4a5SWWNVmWxOlzzvF0qWkYpdg0cbAiVGK
mlNYc9yDJksvJGEvS+vBsWUiNuNGVYUCL9Ey8GsggwVbVRrIt4Hj8/ZnsB9t/tTk
1G7PhnBRiK6zro2GtputMR87mMdetpmlVI/h1Vpb3l6UwUE6YEn/M0B26sE1/Flr
JORGdM3PBFxW9OA5GsAxOXkbQeJaHAj1FvEJI7mukoQWoYywasOLXX5OZxTwMXDg
5MUjkGHMved5XSfaLvLa8r5JfA16OFgCHpwVrh7jabXi10XDVJbCMYIh4habxC34
KvWuoMHcwJ+WNZXaUQJF3EL3+RgmknOV50g4xpP+WsqxED92jxrFseBSJ+/MunP1
EjRC2Le0OLxfkiQ02djXh2KCJ2DClcmnw9/tRI7rGtgccTC2vHmfCiPF1kLg7MWw
GyJPedjmkYGg8vmlNkefi5LaWYFoMx9tt5VScZPXuCeh+dFjdikZkczHM2Gs/6FP
L/bbRsadMVxoJVtdKOvqBe5RctjGCTMZ2O+7enyfNGkG1YLz8YmCwd1LcLLelCZr
5sFME9Af9YfNBcFEv6n/uME8jcB6/c6WQC6zgJvuxwuOd7XnptLbxxsHNZWPOWni
R7LDrxg15Ay7Q2k/0spQGeFO2aH222FRKDTahWGbgq1j/wsiNFY5dKNFH/xfK9jk
5f5YHZ5Vl9hoUNYoSt8b+myvwPjs++jNN8pnbsAXaNaadIv7J6v8tcQIJ2bDFt2E
4pzBpjQC903sxvaMlCWagTgkCwsXZPi5GJm6+FkyKuBYA+Tr7II6tPOYjU2zMRct
QzEIcHWCCf0DrBZ2b1avSujOlZU01H0G55qfDMA18bJSpuMaZ9ANuaT5yKcAqyTM
7fQkYYwarJu+PdZpx/7Ni3PWcf7SWv+KgK5+oRLmLvCJ2e7D8pWYb3AIqy/zS//r
uXNg2OR0z5jxBbsJSBMZk125fsfkua5FehAvSz+3Pcivk0nf+J2ETI2hYfU32lrc
g7LWfejOPpjazi+dc+PI2b8w8vCtu4e7kyYwOjECxifyN6vAYG1OKpR3RDqEt4ox
8J+I2fvijU670yh3++zRrPTqZH2MxkWtbHDY4QJTT8CzZikQbd7+Pfee9+YNubO4
+dKrINVxU7Tb9ePleIGYeHCKm7cHqnC0gqVoszuKxrMiLvD0231pGCzBO7NfcJVh
VA1nNx0qJqn3KFo9gI4VhRRawsdv5+CWsQB7uabCvNixgJUo6wLo+dqELDMqZ4hk
pMgjP63/iqIqmEC+qL6HZRNCQwvrBjrNDPM5Jf30W29brXP+DaIokdNfPdnNG8/g
bflLL3WZtvA/aDBYVMJDLF4E8WhrNxgH+Sjni/aUfeQ1OFArce3w/T1dm+f8Vw3t
WmMZ+ehbu3jCyBW6txHQ0azFHG1rgigzOLhrDCgfYsI8V7uUN40TlwlWDNgyM0C7
ZuFevp6Ehm4BigHEaVktaSHNAHSW4nuruIrWFU++ZrQJpb1+niza2eIcdpdqfR99
qlyubARZ7gqbnItvmRpbW4UpUv+4bnv5AMClsqc/CIAoFGMgitHX5UujPUBJscX6
r6b0gAjOW/Hr8PN7DPrfZE1iE7/X0xco/04wlkFwFxawtbIP/DG6UYzOXuE1XquZ
K9oaFo+xBKgsp3j7iQNBgLjkN5VVGmWE35KTmqy/LYWg/ndwyVCUoQMb2NBHzKY7
PIDjm80ro9+ymddcxFc74CC5NHC1PJifBkMERRawQPZuBFBGSA7IeKLk2ZDcSMXR
NqNlRSXJ504+gg/sauremzyPlzw369J9vYtYjACVp81zy2vChPwbj6bMeXSdTyJh
8kZbdunzSoYqwQpBSo3Qnh/EeF06ui3tK79d9ePw0qtQODaNxb40iiZ1oQ5Oz71/
RZ3cHXuq+p4pFespK688XZi5ygnJL9mqWD9SL20PvY9wTks4BB5D6MuKuEO9rAiS
NWT596K9Ya3/QUJYZNjvEpz8aKViXWafzh6tvDXCkKNVD+2b2tnNtK5/GAVQzVtB
dK/jY+Q/XPhqrKsdN3EdWawTQBPnT5NyzWnw8Lan6sRV2ngO8474WLt6cjnpfKLK
mBKVGLatZlBpx1WoN9CUbGnS8is9Vxvrn2BSE19WLNNTaEwZ1mkiFAxIExHlWL9q
VsY2hHyZZiar0u4r+OrtrrBuvh4ogr7cO+2aX/MEySrc4KpkvTblgUfyJst7nJNW
2aolcp3vXVYa+jihg5k3HljI1wE+7WW0zhHxSpnRmLDEpo/G9RWFMmTEnpYa9qQg
A2tDk5garfIj8pFc9661C1HHG6c+i4bU9toxYyQyXqSAJ8MIBi9TB3Cvyhj1V676
Ast5z/fum9Tr/EABsbf3X39DJfrfgAEGOwVae70FlH4AVpuFs9rvCSjV9ZuVUeIM
nEugZn0SKH45nhZ9A73XzC3D0GpDepcICU4JpxojoQaSGz/OCPNWmo9hj7iUIz5b
yu7l6o0LBfwBJ29RYBbKzNtQfX1yt9V22I05CQPH2Wm/23K/+6StsRt8NYRYVdme
x34cuTPLBeWZH9X6PEi8tER+iIpsjE0P0/UyS+5Qj6QelDWfbUz830kDLQPGenRr
OOxzgWV0n4tVGrWv8hfovm97nY46Zl2h8iwXre7w7u2ILz2IscJSm0N/gvDugteI
1+60uykwjEbqLelF18HZHWMFKzdTJ8gYJC3I0DNnPxDpCQuV11krpLkRTghRMbBZ
XD6pELeCE3UFTVFQwRAtha6ETgu+nReu4rRZxrKo/ikzBl8mD56hhsG09yKX2JVb
KyRCIrojw80aH7e4GaDnj1V/pwXQVez0IZvSkSdBd9GtQyY31+2GM4TsstSIKjiL
PZDmdYp9nSPIKfTZtfaLuSaWe7a3o8wG9NBHBl2TMuFV7v1wOpjOkwFdwlS/cLLr
TKpHlkfVw+CRcNxQVbqEPXDvR4D18wudJJz4umYJ53C36pf5cADIbz8xXb3OmbJj
tiksO++Jw5GeqrDBKaHYUfTaEfm8dA84RV7ABmQJxwtYPPZbzjPNpB5pjSnrgQza
k+l9LJuXJsc76+OUmq7DbDt5jpj5ohrfG6cBrxHaLa0fIxstlo6kQC7Gxm2a34jJ
9u+hMOiwnScWMc5OrjBhl8oe7QN2EU/qu8BagO5fvEkRRv2cFnbIRHbGTOiMpwl/
0nP5fyohYIjsblvYowg0CHpfHQ/KCjPa56ayOkovVKcxjR/ri+fdCoqnJYmBS5NV
1M57sNp5HcEc+/R+Pk6mbBfd6uE4IWYs9YLxp16zisu5TbyMYYCYLOcBnOvhaK2O
T4BAYb9ln3QACVjTLk1MMo3og7Et/NR7Rad34pkXuzIVPKQhZfIxoquHEjT2s5he
8YgVb8S7Ll0ajx8T8aozH2iVt5o5z8pSeKPK+fGEXNPgvBuDcNJkbTYPTzjbq6Lw
u0zmUXHWGiFNd06iOC/Xdsnz23n2wTVn+mAa8ffCS+iznzMjJiN4H2fAbeqvYPQP
pwPgmsUD4/ilhzN9UbshTuwdbs1NS3H8uOiT4WUhbKxuF/7m912+SlSMdlsWA5Qw
lPIiZMdrsr6u6h6BPCiDRdIjAhfzTOTM0HMJjNnwMkTc6zWI62yboGJEDvtahWsb
W17JEPblNptSwu3Fm1lkbZSxrlKZhyvJI1CjXOWuzlkUIiaaqf/F/0NmLZp510Zd
3SdfZYu4635dLbqLkrFAGgf9TPSAVPHanJiiLY1t72qSg9Pyt1NppreMf8ffxbeA
JWOFf0T5khxC0OeFJJEfw8mGjqBDWus/YUk8P5vdQgvY/BYVZnDi9g0VMAeshEak
Llcuc1z5S7RJ/EiMzCpb5sMgWHbAwXzNoG000M5GdSIyT1DeYqw82Lap2kCEzLDy
ndNrjgX/0/1C8mGVAyg5bpEfLGk5rEcriNI2O34UZ/nfGtWMmULRbenx3+6u7x77
DM+0h7eO/YgPqVjG8EwrhyQouHvoUIG8WtKS5Iu8FtA6mFMaoW+zEfiLVDn6c3jQ
4zNv1+Zaim2jh6FYHujFZt0PWraZxqV/efAqmX74BA4MLm9IhUhK8qhOctH8xnXH
8vdHmZ2RrApO9rUdVGryhwrhLE429yufLVibTKdFb4fa0r6mlzg2jYUJ9ixTuluF
0qTD6G94zmRmz3T7IBpQpBZUBRBeJky9IAf3gmjyUyB3FNrjYoj+b8YuzVkt5evq
x6YFZ+J2r1Z2HeyECEJuljZHT5pzVelhkjK6Pw2w44QIZytw9U5tYrLV3U9iumFg
F2wngFjGOUUgCQUGe3R0Ynr2NnWGTtCaX7lH/9HtvZptP6pWjlItxY5INfLMbzzz
WpFh7GnYspwc+/JaDHiBZhuqdQUhUklAROWz0UyjHQwnIktueYkllG6ZnTsGQTW9
zMd5z5R4KXDdRR2UgX6L2oq8i3FpZrePL47PyXP0+Pw4n9dG38KOdwlhokSdbvHm
vAfxRXcrMZGeqYAee9WkangbCWlwp6zQzM5YleZ1Qg12FrKL4WtmjQdYu+Kp7vDt
kbLZEdfEOFheU2EYRrrAhEK8W17eglIBBhLOZ/pQgLGivVSQBByKlRHyuEOkany4
XPwfWSV+qgaKHk+LP36zYGsdFMD9QbOd1tSDqA+KO3q480KbTP81ObfCqS3ekAmM
3BRfLcYuwdFFIFwY9Tjm1AHNoK1X5LG7RspvHKO8Uej27q8qp+cnhzR53gs51a++
oJLuyKfUlGPLllvHxyALoTxFt/5kHUIzgMkPmXK+7xSj5MtHzxO366jswknOIdar
f5Cx5qXiYkHKYOVZPT4CTsj/rZ+4E3JvSXtNrrFyoEisSyFa1rcsT5O5eZsgpF3l
KMUVdK67BaJO0cafIdSW3tiuySao4hs0IzF5i8pQ8DxHZSnIiDQ/DCpk+TEJkAro
gcUIWmu352Oj7J7S61XRkv6miRVWlgpwhyiP9bi/bMgie/Cr7pjl4o0REH04OKV9
5WOvOi8S51a0pXh0G6X2kS6ZGY/rlcV7vHIInZODTAyc6K1FycdTKzOjYKOAlRre
iJI1oc9/a+VDpB4KtnMTC6d144IvtLQPyqCpqnx8IXMZqm3cqfOUAHhLCfhyY7FU
LvKSkLNXL43YDHCUJRSyAUh6R44OEUA5pMGmbhCqFDRl7PORv+9OqthI+XOBHR0U
2joym7nK5giiGF5BcBqFS0C6gc0Bzlv3vse+s7B01gqWXZfFELA0YQf2xD33j5Lx
FtmcCQiJOYSy+U5Z5d6FrXUYygSOdFEtRHw/ygBnpswfthYaeZrOqhRj7UNCnP+g
Ho/QyRpp5uxSM2sDXfX5jRvYyRYVfh/jOm4UxCcW4siuW2HX12gqTa9l5N3Zyln1
a7RouSDgrmTstIeItFk1uUS1cSzinjM6m+Njha9LyWSRv1Fl04bhuDSDPLQ/EFPa
L/uJ7D6tVQfBEHsjbslONEiaZbqXRxyHexYSu8ye3Z9N8zxv7FV71glynzN33+Qg
T12gpMeFyGRz/DAnVZ1sSFOMe9uJtcnGFj9LNP9HMMgB9zzzJY5EqlCqaupsUuLX
4llddxE0KBlAX7FqGEGjeivcMiKi3lbj7B/D/TIllnzSe6XykigCBhKMBPt9Var6
oufWqMymvGtyoHpUDdRjPr0L9AJ8z/B5yW3i/YvVb57g29FgexkUr8J5Yykk5Vp7
8Du6TL19Uq+fwSR1cqBoWqJlql9xAqX/sJrbEgNTGECesuV97ipfM1FcJ4la//g7
MNHhuH2wkI11HaM+57PdI6kBIBUP2oBVEj3ofw9QsApRqYJ+RYr08CTR8uPfHgCK
A0gA7MSKF3wsgod1UNvOpah1PNxU9RPDXqJpHlodn0IDOAEHJILndWtFXs8eIPN0
3zfFEpxIJxtqOJ2n5TAGsMNlW5v7hyJ18ChN/tThe2/Yz8QbrwswLvUgbtrZuWxP
RBbuC2KOghIiBKIP3nlUz4fql1xLmQfbI1trc/8EXGYXIDwdPqaJ+MD7ttUtc0Bj
H5h1Prbt09Fgo9YhnnfoD5a+EkOnmJrWuC1B9MYFJvcZjBr82TDD0qWG5F05We4O
7NU1UUHx2noZ63kzYgfb2sXn6yPRDEiEaqrdEhrq5eazuNwyxzOaNfwRr50VLoPJ
bfKJ3dbn1jP3gYODzCClnB2noyiZ7qH6dksytFb0NaAdmoJo8uacHPICFg8HqjJF
92Lvd1+JeQZuU9XUXbl0731GqYSNghUbmssI2ZeJLmovJ1rP5QTJ+jUa9jPXRgOX
hIdW3RI9IPT4jF8+7CixSx7t94fWNZ5zodxmyQyuNsy78dFH3QUDPiHAc5qb4ZRb
JsDef6WfhJ22t64nxnoeTWS8mJlTVSlNxqjEjG62MxTMY7YlRleG9siWvcObokEU
FjFdprNWHRCHQyxtkvhGBZYtrvfC/o6aVy4QIeakbRQ85LJtEVCWNSzFXstufMJk
+WjQPX28WTT4nPXcHgFQIbI5F7HQKIhaKELQF3wK+FeFa55kEFbm4PIfbJGLAIAt
W0CUFroprePIGvEbr/7w1rVSo4Ouo0rXzm8NM64vmw24WgbUZu6JL4AfXglm7bAA
qdFMcEmTTWvOXzoXNQ9Si2vBFscMysnc3z30Obreg7+qL74wLDWHma5ZzIlyaT5W
vfkKg1XaycP5TOf/RRwO4sK4glPH1Py+92o0dsQZX12JahJNf2FNCNU89kHlIob/
PmqKf0bw1jjD2cKsEhqRxltoJr0MWo+pK0QBKUe2/V8vEmLkr4yWBe0MN7J1BFlE
4NO+zOzlL0rxHcnDrObdxGcXaMGOhBS+lH5szb/T5MmgWBlaur8l9gr0CiF54zAS
JnEa2wEfh3D8s8bS7M+D1BdWlnDfhkdVNSFfmCmQ/e92UF+cvs5gExhLno6/TzK2
CcO9r5LTUXclHkdrWwaJe5OfFzKYNAL3n9s7L0OrQzT7XNGzWu0xkBbCwfxn52pK
Vopafxkbw1MCFmEJnXmIRfLkAw5GxHSDaJClD6nWR+oWHmR/oytl/CSe2tSjeE8L
P/L9fTJLNUSI9mg4RVfK2KcA6sUdfiXUbDLJCxPEIbq0kQVpwLYc5RCqxqr7/th4
+g05YK48fDgwytRRy26z7hBzyEkwlgc66FX8MH33nAOCu410HtLE+vOO9mK1eWHQ
Pv7loeE3CpUXGV3IUAoF5j4AWila9K5yGhdqSskQjWnU4BU7mVh4uR4dqsVaZuhN
HErECHIMaXy1mDiU0m9SB03VKWKZMy6hIBIaZnGjXzEEylKO9IPgRSdHLAnDa3N6
slFBUEwdd2haW13R0uPR5rExvxmac0tgTGMBMogaSK5v4q6OJw7ijyi0P+LK2sz/
V/8qrWs8n4AfmZ8ggdmigt0TcUGEkQ0TvQEuzGHML4P60p/e909kHYqLKOG7HuIU
vJ7rG8C3dibCCT8COnfZl5Mmr4+jSFVjmBKIjsXt6FIXa88bhMy4mppSTqsNZxmp
/jMP4AQLWA36ev9NZ4pY3bKHywIrRu3uqHzkHQTuPcUtJJkAZAlK0IXaEl7/8/Gp
n9e8CIukuVa6me0FxHXc0Pi5IsTq6p79Efnv+g49UWzMKr15nX3mFw1kYksEH7Pl
hBTgzHA7xkpLfoefNx4t4OqJhHCswbhSlR4HZezAJSob1+StlGwTOnn03DENaIAu
yeQKY7E4EvsPczUXRSy+jij0N13i26hdxFQRXA+yCLCKPWvfjj3BO1hCwGFpBeGB
8Ll4PWn7OXx/n634IluNq3k71gdbESGR4vBYmczcJz28Kk/TfHrsMs9kzMY3jyqZ
eHIaysnwOsbK+QiWwEW2G6l+67qVQb6UKzyLoifFSN3rTju76xXf76qGsydmpypl
o7M0xFoKs1yOx0032FvevNWCEHQk6DFxrYrcb9ImcCa3RXHB/XSJfPPq0kWgBRSQ
vF1bDDtU5DqsHQYecbN/FXnXjTszVmByRGxOnJR933NCW1LY5qcDtjZYMWaIzx22
AMIuS6Tpcsbb35Y/UcEryXbzh7WR1zxXDARXkInebpSK7AHnjwLsIivL3vhKWkbj
Ca6di6dZE4lF0M6DOs0bYmbQBRx7lGCn/Z7MlWjYx4UiE4lBT9KFxF/WiiWg/nyn
t0zNoFHuL5+45UCAfP/Rq5kEjUZIXN6knV2jzNOUTi5myuFCnD5THCkXO0FevtVv
4aTlZA0tO6iWaMx1XVrnkW0ym5xiXepfvjOsd6TTae34OZzzTlhRuX481wly+okC
G01rBxqAi4R5lkmNFswfpRvDL5iHd2k+7Bb7WRqz4CU5wXVQw+KtamTvBOvS3QLP
ONq8s8mNTaBp4rwA3qv/AxRx2VUKsnxZMv/IlCr76tNimTjddPyJk+JPdIWFBvmi
/6DCLRUHhBUCRsIW0JQt5NTXd6dfjoYL7y4X0v+F9VHKyY4TDW6wWXJYnlSJ4YhM
gPsaRj5Lyqh3C5nRyTqSujO5IWDE+vtKUo7UD021+xqz3hTSNwvOHxymertghCpw
WMh4c2nNrMZSDQuLE/knmKgwumGY/IzkkZGyTett+k8t84priKzUYpZMU4CCPjkQ
ciPZUNousep30YuaJkalcEb6OUxPI+zkLVpx8ZQ964LEFMatrRKhYm6Ygs82shWI
wvgrcP5JD8zXRYAzaTHTgzBqCudKjWYwdLj8wU/CHuarbTerbLw7GOvtkZOBveit
+BEQfmZ93qO9TkZwwKX4yfIPRCk925/7IFOkkEtjqgJ3fxV9o/d46hQlxB3aQDMF
V2XRYHyg8B00OEnFTjEtS0sb9QAIMVOMwZDMlieHEQsKT9/GYHwV2KXB2yr0oTw8
3ATD/2dTHxS1K3I+ZnCQ7Km9B5UyR8gY/zp/4BO3EviRjAdNAM9xWX52y62WKfib
/8M6z2Db8VOOzQ11uitg+qYpthTr9g19NXfXIrlOpEcKyLeJ6fJEEoE6XN6H9gZK
uDOPwYQtB5pgdJjZoAhCEQ3pZOmHiYcIurWLpz8E9R1ImSpElSDMQoRJLGqR3f1Z
3dwk45yTChQfSr2RbVzCkm5aVgYCgHaIlnYuTxnNDQ0MG/jAoY+z0rvLN9jEJDJW
8meVhDhWDAazX8dGTbzGdth8531fVHCg+1bAC4MJu1eF/RwemLQNBay/9WeYfUSf
l8RyP7WrKLO2DluxvnHMYz5J7dRUTCTyxcHz5oCdUyVvwSCFmsSeVe78jvGMK3O8
FlDfIZ+mlPztjWpkBkJhBiEYBY0syEt1VbsTUPX2zlQwvAhBO9Kxr01hICWmZY7Q
53HGMyjCNZ5UkuDJqdzztf3oRTkubnngIPS6vggzDXHtRjXsG9UDZH5QWamV8JfX
p6ul8HoaUplH5wL6L4pqhOemaJmO9JLNmxnT7H6drvFA+MMO9LjOimy7FtcsRzcB
VCiFGt7Ms81Io+O07fXHQMwEaju7/8OO+sIiioPvIG/GvC78AbyLsskjA1VXom5D
v63uZm6JWB0qaPGf/XZB0/x+FbDfsnRS8yC02ageTt2ihUHREMzT731FgD6PP5gE
p2uIRDv9mmc2ZCNrdMsQXkWqceedNE3qRmmgaLnag0ZslucziSEEd1CEq3YEW727
Nbv9T/ai2C73QdqGs8WJkZtDtREuWvgt9lP7davfZFF1bNzeczSeunw8mfuopYWy
BkuzYz9y49p25UcQOtYGNl9JuzPxtdFdJ29wp7JHgeIpaetBmbufcmwsIVaqsqPx
vvap+oJdoEHxKIe3huNMmYfui73+ZAi41mR+Thrpffe6kgZeplyxoHAdFeERkKtx
RO/mAsMyl+Ojwd0JNmA9ahfq2Yn7WXQNGvM3R0YPmFqR7PVc/HiogYh0gfm96yuR
TMz0FBp/r4JMcljCrxp6u822v4EcZrSSb3SNCaTkkHEEz2jBq2tfCIxqHxKax5tU
duD/iTdaoBsn/kv3QmRdLvnBGDv348OMJul86pebOmNm0UiFk2hABg/jcqvtXitA
VJXDpVwXY1XrNLL8/RLmj+Cpc1Cqo9c2EaBAsgZ/KoFXQ0XQaKG1MMJtMgksCWQT
lHqAHfMwJcbgKpAc409rHSanTccie0vCn0SsidUyze6pJg2Opr/ifyxgR5/id4sT
kUnvb3s6iWc2uImouvTOk7VKUGb8nws1R5KfIBVYjo7rhE/v0dVdGCD+xBMwsCsT
ogPsSrRzZlNpKhwI+TNLyPEpOu/xHKy6H7EYPqkcNlRptMYj9g07V9/d2mWBGFap
+MwLHofY+gtdXoewksEhNCuX/VQR7zMvfGRYzM67oKbWvHdsE9g1g58Ej8OnZLS0
bb7R2EK8ONQ5tTy9I8p5YBhzk/VgFFi6thEZso1oFHNiM59BzI8Qk2ljl0IaO/p8
OsfpPsJMnyHMWlX1k31p5tzUVfBMOc8khokmAqpIhh8xjMQ39IC2Y0z+gnEKoai5
Y17CWASwvOhNV6Idja/NTLSRvzqywe6dAD2HoH411TVSA8nbH/OHrtutUnpWPVrR
IkORstsNcV6o4MtbMoC0wPJss79Ux1wOTi4pr5bjmUVR9zg8OcntiBS1C3rlDF+y
DWOBdl2Y1RXZGhG19wIbJrzEIlW8fLy0/gEn+6xUD5lK/nf6HadNvb0XO3WjjapN
vc2UzcG5UPXzslp67k0grFI+sgtBxU5OtytR3PWxD1z3j8E9LnUIVi8eivd92nUB
ierZSJN6hw8yI0Bj4E2YFsQCKwIC6hb350CRLErPy6Tlw2fKe5oqDBJyxPcjYNRD
1inOa9bFYVvLCJ3ihsnC6RvKlAFgIYAu0sDaL7YYUNcultGc2k2Y0j6Xz2R1t2Up
h2HnRdtIztSUg7o9B+zjdFzb5DG2NIx4UQTFD4r6YstzfG1KXV7RwkqL19/M4eZz
VAhinWIPe5/clRCyVp1Wufd1v/sCQnWJaUXrGg4jKzEjH9W8JPC2DR/9p+kE1CjN
qZiLhVk27EspxFSlnLg+lnE41zoWWDs4+Tzixw7QvCGx4wJ8PD3NoF92esNNjamL
Ia8JKZLvMhGgrnPDg4kcnM/L/X4Z9/yRvFfD3bnTwECAyB1fWuJly5XXwfOrgjxy
vkp4KzpkfulwnK9h18AF+q3NhQ5S+BPnVoSq36qduCzd2NK7Y9/byKuYy1mTqxjw
0fpdQBRdNpHc16z4l3A1HMXzq91Q06pCtxjkNnQ9WFrxYzEu6E3jjChGvUIEIgOZ
ZwXZq636Mij3xviWs8RmkTAocbNFUE62L0iiohia78XozIjA0hcWEgX5IPHDRhIr
kupxbI0QKNTEjrHvInPW2BK+Fhrowy/sxzAcmQwam3iaKYBL/7zKUZiT+u/v/smU
1Sftsl4uWR5d+NRFplUxMrJ6Z6lUih8XEoVQV8F+1Jag/j7hSSoeXfIBLFaEYgqm
Fqdvxg1fCTkFte1I8K5cO3VaoInFQ6QOMhbpf0iwhkg9hYVzz1earSokg/CsJe+Z
W5JmlivGj0JyFzNtbQBeHtnXpqitrnVNkmFymPQFJE9bW3A/1YbaX918ckYB13M8
CK95xvbqJbYJGAyMLFizfe1OGqnMTz89yPBOh0lpPT9n5aZYYhyhacFeS96h1nck
22BfiCfqGGtyMCSLW67T+AypnIfz2qt4mnKFKJjrC1sMZjp54tdoVPwet6cOOi+8
oHHcL01WDVNnTnnz/kpc6Z8ucUhh63JQrNHR22rjHyK2j5jRfcu6beaoDX8qiX0q
7M07swfoWzJLt6KxfjcL58dqijYWQCFeXxuGOctz8fRbZRxe0M96CNDDpXZTLs5W
X34yaieEycjqGYNxtYRztA2O9mop9YTF04GOfi0eTPnt4AnmGscLrFXS5b42WFFX
L2z41md/q8LuqBDClO6wjm9covkdNEAqNOYU+7BGbRLOUwzxfEuOK5zWdEhDBeqg
w7GW9Z11E7hANhwSHYjUslhj1CS/vpMqXPBecrkj0PnEjGbLFTbozZrSTP4kDGql
yHGjYwAgv/RZ9FTUikE4R0S1IYfwETdj4A6rb9OKL+HHNrUaVxtruv7qf89IQ/gt
vwd9kASNA5ttPI/qlyAZruKYy5qAovd83iNTy1eCUCXK4MpnWlJaJF40Qk5ly9Vm
A4It1hLjfwBzhIhe+haX5EjYuw4eQMS+dkCGpaqaZjvowKrPJPLln2frPDPd1eNN
8uBWyPEIZ/xtXkJkzXAHeHQBzMqHaHy5IUN+MetPEFc0TCuCXIpjhZvdqdQmBvgA
Fkpv0FYRdyBxjp+Mca6wIZ9AsHqEdkrF8fWsGxAFwjLHsWy2Z3sWGFEW2U7I48Mp
RbVylvta7alWilXsrgLW7KOsAhDpk+zQixA5C2VeAM/xm5/drKlXAvDAD2OAx0RD
4Li/Q3DiO0F5s5OI39EShKclG8Y1//gLhCY59ovwiY4B/Kenm8ZanjJ27lXxrmU0
SvIT+61FAeKk9tRxTiQ6k7ZldVUViN6Nw0UTiQSxpQJxw1IpiumyFkNBwz175oBZ
tl2aiPtEK6EODNwaemBm6JdM0/HHH+thtaTeo8zmkCM1a+ee3xJrgYkFV6/hYaS4
QxF3aIaNvZo4PkM8/5Cv7e0XhRz1pG9Ze4h1LNp3CbEi7bZI/qFkoMvfxCxNeLOR
xUqTRAqOWg6P1qrzYFIBuCSf3y9OZ2RkGFpXudwD2cxNnsnZW247lInUzKLrvhwJ
ayBgrBjLoHDLO9PaFbGTBdD/evx3ysqxjyKEtaLDyj8V1TmNG7NU75HwlYRC7yha
fUrWtA+WFFMbBVvQl9EGIhdQDEHMsfAwfrsaFPM6P1z4EfkpH33a+pgfR0MkMb6l
Yevf4DH/lYB/l10/IfRYv+wlj2xSozY7qQ1xKkK+6HZlpUM+2vJFlSuJ5QMMXyhp
yEF58x0dVGqaHHSTlVvYWWepKQVyG4LEloM3FXTZqrn4cfgjlADYm8JnC4bccbz9
3twk9Tx6B7Sgqx3wm4NU2cKcx/WdLB96SWhtVXt3qEYjAaJ06DC7ZrlV1ePgSF+y
LwIcHJ3RS9idae4QdfFSgj/YmF37KTwvbvId0qsH/3Tr98kDGYmTYvZ4edcr6wg4
9Px2e3oCCpcZ7GvoVIFsHqSsXZ0lXNubRXsplpvcllkV/tTfj5qYwbCms/6CLfDw
cHfeLu9mwLV8amDVnJxe20eemjlKScbGFaVGNLUpxmR17pgINv2fWkVhnAV6fhVE
pgpWK8LHeVCkEZolgHrHmbBx/fUja6+GmZGd7U7RefUPw1pK8sDFLMFn3dO5lIrh
0FszOkEf8OYsiGsqjvT+uru1W7vwLNFKeCc1RNzYIjuC1S10UZ2YzspUEqbbFmUe
BdnQLgiSSjuNXzoQSVZT7Gpwy3hP4abC4eMDHBVoaI2LMQowJnakQCn5yoY9nTFZ
VocAIMpdhhSXXSXWZ3maFGtPRt9XU0S1PF/VDVigx1RBHcFly+LBeDKJ2H3rvHhJ
/Pk1rLnGJJMJvlNs4DjLRwiGGpHRbpSD7NSHKShe3zHpmfLZlv71dM0DWZJ7vCcq
lvAY8hJRT+QuxOGiytMiC1PQy806R5hEl0bWFAu52+YLfmjS4xvdLVoeC8yWh53y
tNACku4lWhS0AWEP4LrFJCykdUmHowbfgyi8/F7LV1h3gkUo64PI18oc0XnGSdii
RJrW5AdYNP/gRfYKqr2XY1Zxs28Vvl9FaKpGI645JZvIhJoDIJjfqM+YpdioDFDa
G/7Mr9gChoY3j8t0q4rL/FADc/jMlVxkuX70YQDcPlCcUZjFgUc6u9kuM8nQPvRm
gcGYmJPG1xPwW9wJaYu/4dSfOd05D15Abg3vwfsRJbE7i9KRrsXvVr/QzkVp4o61
sf0MY0xW2iL9+JvSnShCL0QpMxTDGaxf4LuSQBbdZ5ea+E2DMH3FhqCffHAy3Srh
x3cusan6iK/rqaoU0UtvA7enticz37uu5ghZFxHnjniV7ZC4w6VIwIXwymXUOvsQ
X8tX6yZW/l0HcMacunEWZmBiie6tWVtjlfNAJR9ePQ3ZvNxMbRUWFwCBWq18ijeg
ktp7YgWC/W01N04HiIlemvUE8Kh0pDujSyF3pw+8sFxIN8KnrHe/3n+Hr1UqG6md
RfI7MMhNSrCkirFuH4Dd48PzYsYR1dVO991eNG+udix3vyhRUYPiKuK3lZ9JRvay
/C6u7vLX+kONorzoHWpExIrvgZoh6Xmq68E1asGa3R//XFntDZ73IIxSuikcVhch
7es/yX1Yk9xjtKIIbCdXProieVVwHQLh7XOu0XDBUCr7JaWurQhQqsiex9gz0Ruq
Z4daPJH9aDyHNnkaHv0qc0OaE9I84yiOyHYtSOYyWVQLjH8giK7XURW5CrgL9nQN
8Bg7F+1NutkTvpjRqsRaYr+Jg0pkuxLNC/Lf1MEveSDK7QdsKvhQ3gUIODFfrRXZ
jaltCu1CocWv21PXvCGhjiQ47vL1ST+I4mDMymt/hMgEoKhquOmDQTeMP5Nw2qH1
o3YRufisdEpLaM3mGAuJLvhMFoSvlu/OhFOZJNxf4sDvq21llPMcB8GcNCYs8clf
ajEDQOZCi0jlhxUmjR6FiBA18DdbQzkfQ3uDQokW78hQiFH49tWaB0TAk3JeCQ77
ucN30zXl1/KOFLqkLi6PoOKnItaqxQHaiKdGW0UAknyYnwY+0RLBLN3UPzg0KX+i
rgyH5t3ZvdJgEkPAi434foUexETcCK9MuL7s9UIecPGp1KOnTBZQcdkiaQNfOxPO
tN+/cgkGFe/Br8Zq/lEHrkFdJcvu7XVmD5y7DRl//m5q4OeurYNoWegmwFZsPtN9
qE+/d/+o3dP3QqZjcQaLli+haCqHGlBVGcyJfCso9Tl/Bo4FB9Xoi3YpNbAQX5eH
UhTCnUMenqQN6bxE4K3DJH6gBTlsd32hHd/4IMiot8scLwSYMtDpNf5UzoSBsO4M
rSOqV4krFV/iRLkdStIaKs44UYHBJpMEHvPJkJTOB46MZfTaWQFQQ2eS5KHF2QeW
AiwIYwBGkDMhXeomkfNDguHQ7+Ow17slfMWuDeElti1pC5SUjI3kntBlK3eX/SXB
013Fp8PfyCGW9jh7yTTSuuVXdKSRlAZUd1i27kFWYYiWQ0GhAoBu5YmQdln7hazd
Tz/yokwx0+ZLGe3URXvgiUVltx9b41ExDUizy62ptHStlBxTaGP8Ejbc1UlKo9rk
33WvuHmR3/xbfOWKGSRCV2/GU2YpKuQjPW/XjttGBTC/6GaNNsXwodm0jedmELTc
M9iCQJWomrv5K7Lm3403LqpUg6SYuECah+M/M4jbqNtjZhi3p0/J1KFjUIUzYa3B
IJvXGZza1U3nuOZkD66RyW1S66HvVftqlaw+F07lNVeLdVOLoweypiz0kcl3WZvB
24qFnjs/p0TX1eqj51apLawlZPyPX3K9YaoEn2WajiMW/DXed3XsHM/42aZrMQ38
Ani3f4XVi+7ybdBbJBRPHubR3LAvVLK5oTZBNKzks0/cP+zVj/kpvyFTOHmlOG3A
44EyERKPndBBq3/dRkLM2gUuuhrR1VIN2Wg5Uxtaepvkb9wLJOkxzXC6znHE+t++
1NyhsjJRjW+QHknj+pw/NA9Jix2RUG1MwzQc0tg1WBJWGb3NhcTJHVUA1VL/25DA
Y8SXOE5hcD2WW7fp+lhHJ2ZOhaSykZxkzGG2BPElBR+1bxPSTNOuBHuFdVgXJjck
yEW+fn6hZOSatzL/xHDZsfqzMxSTSQUozcPKw3byVmonCDJyY2lJkhtmoGzd5OFn
Llf7/epO0uZj2mSm/hlGSmXS3fWq+bwjlzMQax2K1e0VvH8s7oGiQq3Al40Xa7KA
XdytOag91BVqqtIAAuSzE67vCRHsUBgyJJulZjRf6melMb96YCFXYfSiQo+0nvJE
OirnLaM+s4P47e9PYug+zWfJ4L0S/TO6t20p6OrXhtFRjk55HekkDVLZIO837sdV
tFJyeHk1Kc+RqErFAbGnzNpAxteu6wxY9dSKT21ZNn4XrKVp5w1UT/dW/DvzrLYy
2e4hht9feg6vU3DKAUSkm17YGRJ2BQdIFJi0UTdH09uoIJJ6IB5rXC2Y0y/CkouT
qpr7gFIII1TxXh2tZcCd9mHzP4jm8R6yHe/H6IMCYNEHKtVVvVLJv/q7Szc7/Pxt
4Zr4kvfwSgevP6/lKffzX2nY2IHa/pXILaTK78SvhxF499un0kQJZiZc4Dk5VsU8
fiXmL8IUWyM4pG0WPAdyeGHeYl+Kmm5F384JIuFrH9IG5QaYQEub9Q7omQK/lhbY
bCMNr/y50Gqq1MQEFeAQWTWdWzoLuDQBhGg+Ex4uc7z1cfB8wQZoX7NIkij1pbEv
KmaumZU2Ip6+GpvJqd82yqDuLCmvUYwGJ0YojTmCWlTqUBQ7t/APPUkAITE4shZp
j8XTwoOzuLerEbLU7FywmK0AqFxXc+rY08SrT+hrxkR/U79vAd1fevrmv1OI0dVm
lRlGMhV8ugC+QVZpultGIUfLo42jasksoCSFuuQEcLrvULA4I3iNT5I+YygUc5Kd
/LYEFp53Bgl3R9IKkZXFPLW6K2OzlPkiapAboTog2zUWC+GVnHusIZ+q4/KMQqiO
k48G8naLicPFYa42TqVafC8hTfbmWqq6ONHP15HhQt+mwAuTdu3augVVdRLyqSof
Kt3ahmeiLDWrCxyVyYYdnuaw+pQM3pQ8F0onZiBoXaDBAMXA5Kx4LQmPW2zEda0u
2Uiq2KOiGt6g7Bb2b/ystaOMAeQLgPMDvmxRXDBVjpL+qUb1YXclNtPM5e0Mxxlh
emyISgaTNLYv9BDffZZ1itgvAA4/syY+moM90lqwrdu1ZrtIZFdFHiRV2xEjctAX
c8cTqAtt8j1RhG2YFAXDiYSKiWZ8KNXc57MDfGc+2W9ocYJwQU8xpMPPUGSv8x8J
V/TI5RHZy8Asu1WMHoBPyIbe+5Gg4RzEd8Qcde21RtmOAQI2DdDohP02Qba7Tt9j
0NMrwQ1d0Zih4kt8DnmwzzMP1CJg4nedJmU5Jt/ZVUeDeS2nbY8VVLxtc+8zK2E1
9YccxJ2Qf2wL4MV1iE98y0xuZcoVDFyn6qjvK4cDtU+uwA5QsBlQXxIY9E0CMX3i
/hmrv1dtG9RyPfZVRwhhk885WkYznB7QyDTA4jKKFaAkeT3okXpJeqeCK7OlJoQM
R8o0LxBmIwgFfZwnJSz4qYxt0A/VG41WH8qj4ZA3Gy5CPSeOQSaw79DkN8tWv+cM
sfI6qlUgq2cu9CSBPQbTb4XDSN3MQ7GpZOxhbmIT6Hs8MSpWWyPJCWitVjPvjt8H
FOlwxRRuLJv4pD3oPLK3sP+tkDxKsOo50/opOnDI74QklIj25aXNtr3oT3JsfrIx
tUjwy+hBRhgJb2hci/QeT4reRNEA9HYSUEWdi5tN65XXX60Zw1SeNC/YHFNjswz+
mZqOym+V1M5k+ZkyuIcLTAxxsUbiL12Xv2YBy7nGBmsg9voMtcjzPQOI9SgxzW7Y
BGniozQpPdt3RPn7779KyizSvirkLisq2HFab53R/wLoX8yelVhBkRmv5gY/lNKY
Iuhe1hUG/tWEQNXNYxuM+pyqa9H8gkRH3GGsM1i1zH2Yb52aGqONEf9kMFSC8pUs
0egrGrLqsHdwEcaElb9j6a7+Xm/3SeJTdbarxyTyEtr6VzgG+ATLBrG7dot9ttnr
vQ/32MOczIsazROr9hQiwXrhVSJnCTBiEkm3giqCwn6M8T8jbw67C5ZUrADUtMWx
sj1ui/MhEfghkUGXEQi3WKLTQPRiTBQJNaa8OK0DrHWu+969fZLLKFVryjBN65Te
pickUHsAGbYptRO6enoHjgHe/Fep2fIAhnKwzV+eecwPaGtQZycbw8ATFe6sSSFF
c8gimpm0xFIfzEEV+YvH6C81GBeOCQ1VIJJ2RheltS1b40D5FwEqf9IKuNFw/0pM
fyxc4VuPrKmB1Q5xZGWxG6OLAW9ygkUaoDkPo/fQFKN+gJASFMS1ZF02QBWp7vh5
TBbahlDdlPF9kIteFrYK9AKfDeo83l1/YgHnM7B8tg9BEKTjEU5LBZOEZp0Nv/0W
9PoUlbuzpECM9Q2lIe+f0lmYK3G0obZ7Qu84PqY/59+pC+kkxvSB8x2mtFhDPb2N
gRsGX9fe50lFOUGzlWQx31YyHijd2Tr2GEEILYqhObV4gsZO1xk73yWVpOWH04/D
YoXSL6QrVNCmxDwQuvqDqjY7zkg+53Qi/f9ZsGn0TRS7dwpAzPIN1FUwtcyY3Mlp
ua3EgU4Q5njh/vbrsB1TIkHB4vmVfOYQBLLJW5x6LiVTmMivnX0Zxa0Qx7wNR7s+
nb8Qo2ey95ip36ossQAb0FnfdcemZEbP4uFzuoApVdoNRBMJLs+qXxE8dTksIcEG
3kKKMRxKeWKdSTC7CLYYNlT33enylywKne9w21tLYbXE199rp6v9lhk2PVoBVphB
WUoo28M0yZzbeXwUR0dQ0ADb72xhalZHtvAJMOQGn+4MGJ1K77p/VCnvtGuLnEhN
Fcf3w2tqctYf5LfhV1Pb1JBSt9g6HTnsXyXEdfOIpaQNW+c0CcU7lSEw/3eihCca
KGsobC0BRQ6ghmnh0tbXTh9XMPCZQTo/+t5mNg2ic1gaJB/OO4z253s+qEStqwgq
QAsmaBS2Jbb4tJNBdHNRPYRdrp86KiQP9Up+ugRxsqUwLC6mkXeC23PIHllxQdFu
QFG1AvcVpk1wFkbTK5XgsuM7QXB71fvf+/m7BjOwgA0pOoEBfqpaVW+yL+f3k9QZ
tHr0TmhjKHN8g2DDHX3RyC+azdT0PgDmMoAyZPbOs4HZbQznnAbyrSuuG0T1Ej+y
LXcs7r/lXcSteEkOnmiiK6CHk5L75vZPrVkIc3NaqdpkavhlEcLu2NfzaGPRMB5i
UWnFvvOdFqPjdyfFOE4gNjh20sTSyCa2vliR7KygvAEx57hGQts9OVRGsxrjSl1i
GPnF0K6uQsNCR/p7F3lyPr+ApCcNQnniewRPosumuvpqnHoSPVk5vxqLmefCLRoG
LEiKBl0yGU/XBQJMa82x/aboBaNFQXXCERFt4Wi43DviO9BQvIUV0e94mwl0Eq2h
x1FCei8Ne7YN0ylIXa5Tnu07TPpajRpZDDz3CRaGdeyXbYttNaV+p6GGxYhBoBGX
aslbzovSPdS71nxRiQBwz+jPrzHXFtM48Y6vxHB3hIaH0U/Xz5djL0XrmxSOCC/k
N/QCznjncvc3EX1d2WrImsGkEZp51jwKieeqlfIoYdYn8TVqcS4cvgAgxijV34Bm
onJSXs1vd1//wKWtcfBAaAw/L1/5AWZhyPDU6GYey2Su0MM0QQkSHvcj72RovAGA
XojvussU7iWXEHIsDkzbeH4IrzvaV/srkj2vult2WrICrTO6ZHsZd0uALxFWpqs3
xwaC/lPRm2N3smGtscoeq4B/R/gv8mcn3ZzZ7QwQppLPhfiRD2J1447ofNBtCKGC
1nDE1qgXL5kKYDqiD+OB10zyjxskiayHz+7PDmUhnjP7U1DhbO24UsyON7t6z6xd
IyOcpGWj0KYrnTNrudGuYh0HRpyu4Ge1jGb/2qtS+yIeq9RYUqAajaQNd0yMyqLt
3blHRPYJBgq9cky49OIs6G3CRYdQ82X9+NqPn3DpjDG52f7qnGHTPcm2Arhdg1XY
Hfs+fiL5vkkaxEIOM6buPVsXo3F8MagWoYwiAQD9Q5yb+7/FbixxQAqOqfYovO7g
rj3CO/UeUi4pOWl6J7+wNEhiQtk/IxVZ1bpN0h4HOyOISwgM/gW199qcV75DJ3pr
q6kNYJI4tCcYChF6e5U58DkGr9XRvoYX75wpv0lxbutipPhQYQRZxd8e4LZplwxS
xFZpnNdcs5dAGmN5fmPzjVi+mQcZlnoZA9/XEvVuuzJu/nY560ADdlHp/1vcmFKG
JB2ENA7s85AVFE8Ej4kWsvK1MgiYDW1nW8mHEpNL3PmRKJDt8XtvJL3iZMvN8hk0
jIexC4xteaZ5FuWvJVgHXChutDyu/U6m9H5cBc8yZoCTiEinRgFEYimJyBancCVr
oZlYrXGBqUpgSrh+BLGJ5K5bcaWZzrZYHEokBOq6vRhAfYegIr6fjuxGvyCcTVIA
00zgtih0UqQKbOvCYdxvL+HkSoU+/7QCUFvorTVQzF5q+4RGemZXAfTNGUC6okWx
t1L0nk+CjZcOH06iEtZj1YFa5sfYWYY60Apv+wP6jGr6iOc3w9n28fbWGiXuPM+P
5pALTDsxQsN9C6KK2VZwrYwdYowPs8JUR+6WpfdufUnjNUyhbTmUR0Y7ra7PzJI3
b7SPR+JuzaauEzihuuhh1OgPmwCTL8JmnYkFXJtjfyDybRLKdGyITAaLGRe1nNgd
5+yx8TEC+afJ2SdihiFveua8Cr6vmzJy+oP6VH9b5ssJFBlLf1dtLSEY4AC5VnHB
JA4etvE25Js0ynuo3YPCC6//ECxz7S5uN9DIINzhW28xMUBMKTXfzT1GwOwJXTZa
TrD9pXvEaAoeIzFG2d0oNLm+fYGxGtM86CapJcqeO9V05l6iE2iFmRw63ivaRgkV
/Jv/7FICdfnfcZqvQeDn2kKqb9ZIQmQ9am5otZObqH9jiW9n5CM2M6B/pK9PCZ87
ASi0VsJKpwTHv7klF/fobYd8MWXkR7vLX6qZv3Zs6gSJRLaofSgzSwfbjQNUVdPL
QrkzQWapkg6/TyW52CWSNxxVWS9mNagpEfDahEkRgclt0GorylMDstj7W+ZacP/G
WL2U3lC3b1KAAQhZwuwqg0o71sXBQNvm5W9hI2StO0TgWyTb7ziOppNmlNOEO2K7
A9oaYQYK0JcP0f9WxYndEcWlTKKWirL3jX/Qt7ocB3xM6eulFKy/QVw4x3St0GFI
50heHF5CgoS3GPfMauGdRzaaJD4C8qDBDPTQqDacam/bXDdXmaQVyerFGht+py6P
7QzwrdsU3sVKKqQ41SXNeLGONRGUJPZuXu4gILUOA6BP6pdfrDKNR0nJo8is8jS8
aVRhilmLcK6KhE4bwQzUXWKr4xRBITw31VSxHU3+7ZGjPu+ni5JHg31r1+19qmpv
b4T+1z2GNhW/UmoMxU12xqnPCXgo2pegtzRwHEMQpMj762Xjm3Jo4XWJZReFC58B
hy2LNrMEfCy3VeLvrVTDUyUJoBsHcs5Zrn8oWutkwjDnm+44fV20FqqKfmUxNyvM
ya4OCneaRbA3QRZCY3apV+yH9lzIHZqjk1m1+wKfrICYEvBtTFfzTrGFRQpi9vg9
e1/y7WIqASjZo+mUqPhjzSkwsfoCmv+OYhTWB6+Xcte/NKA87V5C7FBKcvH8K+xs
pwAYK5+5aXkyDkXTYxI3guV9PE/pxR4Rmlht2V+N1U24vQ7vJ/I/4pCnsaEPfBNO
SpACeGlfQRi2JJMQK+IT1ze7Z9zODEvFjA/uGNRxRp6pSql0ZCrc8NVMn6IqIn9N
ahxl+gY6jf0KVS+C5BXHZefUIbrufsKLY38XgpBY0jJU4RgUKWW0aOwISKiilbjf
pKHY0LBYRaw9Z3vTvDtS+k1eClWwhX3pUA6xp/FmT+zbqRZMef55IFGX4f+sj+MD
88SO1gXun10zbxjJKqeGqRAKKsLxYFStwiI76jQaPYLUgmYSCTWD0B97GOv68w1a
FoM6Q+cHOqee+UQ4ExAkRcUjdHydMUqxGFzv9upASPIQRlYn/85uS5uOoMSaqOxJ
EqJ7tpYyTG2NGd9eUFqzh66VVA53AcQvDv6jpK2Ks5y5VCHEraBEKTvvFWjoApBj
vRC5cIMxKn91o1S1fJkkM/0iVyPO+7DdgP240pT7yRz1gxNxgEq2Jd/uVbFhTDVl
IDxBi4aR8wsRdftiamLXpdC4r87gNEiQ+PGV1pqTSgRXYJQmgwoWSL9RGG8INd2Z
AgKfb5Fc62nDWYtG2l4cfmvJkT87RwaNHr6bJOHg+/rSzNSoJ7Suewn3nfHSIINa
vxPXwqBtrMVpLJWps9m6DqqBWnwxqSJrBB1rZsTk41D/hCefRhy0v2KYGmQ8aS/J
q6PBcA81bvF3kldVxaqjuMmAt1dmxmOfaPP/cM2F7XKN2Z+hBxLmZ8zriTDQzzyN
DaIYCIGbE4U1cfFsbm0UNSjuj/5ZWv2c1vfTc8dDJEhPrB9vfZW8g6lOugD58W8a
Gx141sTEd7d6FGLwoeCyGMfGV2ZpHX9GQ+sGr4SyOdJnwK6aQBXb5T8g0wivElBs
m7ZaWgYDFKTejMmUsiSvtx0vMhgkOm0zFtwKHC0R4GXCXZoXF5Z50MWJoCDVyzoU
RXlm3EVYzsYmAbAFSLWmiqcgtgTTVPhC/hcto9RTA6Fy7kvjv8c25jwM4TLrlSL2
R62IXoMdVGYEBPusKa/Cu5S46Sqm1EZ5ZK1qBqgkmYG6+K1AO17Bb1IPkFUBjwyw
aJdU21E86H8/AJXBawNI+1K1ZPwq/qJioY/0TFWKwI0f+swdLuKKQ52sS4pT4C5s
lnYBfOj2qGlBY71d+z6lb1mrQWe2lblgo8dROjwKnntk/JPmrxqm+zFmJyDfWqgp
kgQPWfhlHULbykUYEeumLdeQkd/5srp/+Tk4wCzGagcCXrcaQvx9i05yrUuN3Lwi
uypIUGjyyKSjCI76NO7qoSRntFowJDXgiibjL30PREN8J8GCckE1E4uSws58ESpr
M1K75GdcGV06+qHAULrXm0/XFfBnpd1YJvq5gi8i7iiaMkvW0TWcGfGYt27L2Y9w
qIW1zPhudSHxmx6hqkeIzl3xEKBRwjeP0nAAMYn+fj3yJwPp+8OGsguOU0vQXTgE
rAOHAoDaS5uZj1j5lhiA+sfBgPNzZf0sH2IGIkHf2ozVEqynT1WB/v4elo8/wvZx
YpUdM9t9gSvuNzJVDqvA3jHc1KeR0LFeVIhRehnNbTY7OLL6/BWZGXw1q6LuWhld
AKokS0LxVL6LTYyyUqkoNGJbHT7znNrUdy56uKn9t5XdzL3Bq/5zK0YauisrtwAH
7jpo12gCdNdPvomWcw9DjoXxoLJ2jh2THCg0oYS9zg2316/Li4l6W5MF2KpwNw7O
liqXRDMUgRRL6O/4cDtYfqsJoFEqOBYmV4CsaldilE+J+vnpOwoLZbx6SAFXh+eG
yeM5wtNSIo47th0xAXNV9v+9vzoX+Vf0eApboCiMt3TDO1IMHS1+UbXWQkBT+F+E
MGPUfoJdWksEfSXvMgc65cMSwbTEO1JjK0aNM1JoEpWJucKk3yqc7U+9AelqgEX8
eZULJqoourGAZMr+I555YQss7iBs08LZGV+iZ/K0pP67cE5AnX1knqu0vCaoOqbS
+3CyjGv56LFTVJtjmw8qvwbgxuNejC+82zBrnVbc43kczUZBH7m1yZJ/6aXLt/AU
uFiT1VDHlDUVqGDQ8/hn7r02xX/0dWxxve1dn6miqnmmSb897vQcLavUu+Oo0jsI
VL8Ap39q427WmP5d+bXMsd15WsJmiAH33+oMqIAKYafPgbNPP5Ou+5H+0orjG2hM
DPQaXoAoA6xDqapUo0F2v2g53gxj+5QBFIS5rTdfHygO5+21Ik5xemsCnaggmgva
VVj2yCQLK+IO8eqc5EHqtRttNc7FdY0N+HZINhrHzjEAzrrsrnh4nXB5LOKEuOkt
4dtOIh2bZplqi2HiIwRSJbwBtg7LmaT8IRlEM1xDajzXXEkcce+DeHcagFQQPiCf
2K3E5D6DdAGsB21HCLDtSkEt+EAyFk3k6WdZRrX4jS8Rv1b39ErJvaJYPCGwB5TP
CIW7V7AgZ5fRnJwAW5A1Bnh8GNmFTlSvtEnEj8ul4Sqyqj9WQUYFWemwQ5mj9GQW
OrH7Jrhyu8JkZmiqByYFpq1iuPM1vcK1Kqmb3K0q3ZcBXZah4LqCf63gASet6gvY
b1dMkVRW/8MiWiuq8st7AXyYYj9YGrYdDkCCJUU4+Sq+Bi7Ew89ip2aY3dpTMiI+
YWz/UPYscX7ZI7tTznIQkfEmxGVA5a25ERFHw08cc064TNE6kolLzdUiJ2VUtgIo
kUENIxxx+LEDBFq8IxDwM1V9QMzTEE3RJfFvpb6a9QeP2cfHaLMci6i3LxxxIBnN
w/LxhWmW+LKDehb0cuo9lZ4GFseSVqYQKIgODV1XlmcEa7bRO65x13lAzYqgMN0b
vUm+TH5yUSObYbIY2Nf2+j6CTkaobC/K2madoKxgKYfseK9tcYph4C7Q1EMtTk0F
fZLo4C0lwlkHRj7GVkLTXgycs3nUTWSbE2UEGx15fc6XY9/O0EsVlibyMKJr+bDx
m+qIT7eCQzllbeGr38CaLtMhDMrH0OprYTC4GKtTD0oG0/1OQqeUu3U14v87xzRK
DEQwAsVxb+LjotSvflWrllHRfZSUslkbwmMHYtYpMCHzwfIlR8pJ54x7Mxn9/nI1
xNSl2cl7t8GtAVuzABoOFgOZakAgVjuu3d1kPUl7KAIS0UscSPqCL0+QnmyczZ3o
s9oPv9zPLiq+JUplDVRx8osQiBS3VuhA5XPpr7CKtAI3VDBN28ITAj2oe72+yrWY
L3/Gego9dJXRhch1HCqTin0djL7bNtj9M/UxZONZXcjOMmphKl4GTh/Ukj9tXoG8
hGY4CgYZV/gCqmcMMzZU3tQjBNYbMUgRcdhFMGdwRcgczSF6gvilNTq5nL4etw2S
K0ExUIl3MUh89YnuWt4CtlgoaUapgn9cwJJdcOgDYSaWd1d3OY6kASVgGf2risyT
CKPtg16s4E2X2+3Y/WtBB57JSux47ScyKy+/mTaXEvrw694jmrf46TVVz8ppiMLT
bxDb/3WEHKSB0UQGOCqYrr8RWhM0++DvKdb4z9LsZGM5HrzBbFkVrrzKbNrUMgW3
n8tKgQVI3vcHU5Yo7wErmSaKroNhyitsFuW6B3bbcF+D8AYPrjIZfmrFdK/shns5
v8Yj19PoxajwisPD0zq5nt4bcfjZOGvOwSqFpPcxblJraUypPv5+4KzGM6wVhghM
NjroF72l4GCYFKngyN+EEfdlTb7s8SelCUnux9l0VLjn5IkqGjTBHzXf+XmjVjjU
hQk4QVEjESPQ0ZYi1V9RoX4QDJGlH7piyfsTHA6NnXA6CSy0wr2jj3ctOeEt6/v3
KQIGoNvqQDhQ9okeO4AyarvZ70p0Jo1AkLB2VPck6qjediHFi7a7k0/Zf0mEMDYJ
GH9wTOayTVzzJEHQmd1iykab8sNj2UGrXQpT5iB/5HHMAY99VZnSWMcgMsMAZUzI
jMgBtJQkHeKBYF20FGp9FjN8JLi7ob6blf/5vmx6pnBSATHWIWvvk2+VDfkW2+NX
DfgJXku7AN48Z1qKiREVjDiS98QeT2wsmMuh9GqkfD7eykohPGKIHgpFGnh7pI18
QbmTSTpHQSamLJDOFt8PfxIO6pEeo3DGUj/fOuZY8YloqfNqu55FQJid/p+oFlB/
oXUGJZbnsy37yzQMTw2spv4xo/yHCRUpIfxWnoC1EavKXgBjGJPpZqKfJLeplDJy
uQGk7Si3mQW1QrfSjD4lLvBq1JEY3CjDu8bppllPqVkGdgLACWnCWxvQt0fVt2dL
wxsfX9wl5ygOzU+WULQpVLS1BnWQAcECUQyo7G0dgSGylOY289LAl8ZGHJz92aRJ
2jnQI2NS3H5TAtfYQbHwYMll6ABRSciiCqD+/tsz5oeEeCw0yyoNmL3LmDxzsLO6
7v0+WLjjhnYj6FYoUDkWNGzwv7OtOVvx7fkVuQqX24AfaxpIuPb9X86JpaAVpU7G
8FW+sSBbYt/HuvsZH8kjrlskEWvoRp0fNvOmTKG3h9sxa+IV90ERD5r0bPYCadI8
XZnAPSsDUAK1IJ79HpG3HdJCGM2lRfybePw5S00L6JU94FDii5RMD9R1RK48IBfP
1rnE0cHMZJ20Bi4lcsfc1G3ctJVfgfPe5j0Y19gYRxweU0mtxiu2iqvka0qzcK4K
tewyG+tTmiQgmyQfijhlOLHE9nJ+0nS2s2vliry9TtZ0FVsD47KZoDYs+ZKrvn1t
MDjsCLjafrg7Qpks+nKk0DZcbWfaN5YrtcK5N4p6VU79DkfmaKwbxjcXsb9EsjOo
Bg30FtbP9KWMIo4oecTifYwVa2CFzHt63ymNW0BGw8Hrb8cXpVAgbV3vnFJHC9sl
g0TE1lQLXiM6Ixv0IV/oOrmdFkozAWr/+YCIlIgtDxzjikI7UIoh6IkV201eS6Gt
EkZkiTg8hLgFqYRTw9ZXtSySX44zjCgLS/NDwrpU1MvreDzUnlgeRRuaWSoOat4l
+mttIhRISE1tTw29M+4jn6CA1YniX5vrF6ooz77/bdDt7Q/EfyZ4EvR5GpZio4xE
0xlOiJvG2gQ7G/+8L66MXuxdENm2Ai/73C8ZXtkdJYhBLBudqHUyGNIdVMtc7nQj
UE0cfI5WaLhMQYiBlJZ0pbzjpu3NW2eyMBgm9ZffFP2poxSvMfkl5bsC54VuMlMn
spCCUcd6OJfjGtmJ355MGHigchchGswPtBakbW0Rs+KaaNrgVkIbstzJVED7WkCH
MWJANb8j5oa0wgFXZnSphTprjxyKNpK+t51M8dEZmXCfa1yhLueOfLs2/J+HEAc/
bSeqTdDCHCg1kJTgnLN+fT6U2I1/sLAtTGhzoXF2CiNl+FqEluVcRDNU05jRigxd
tgmB57TNfhU5swdELlLHd4xdnG2rK0WAGskmvlxo8kucy3XhQsGEsiljVhANfmuy
oeRO+RSGDQALhtY3SAbdQgZcD4dFRGmy4O3xQIBvNYbygSvrSS3VAiGacQz6mQx0
vazwL/MEPI+tjH2T8wX0thLsP4/XXEZfpfeSuFVrxSg6ulJFmACTKFUQs6wdvqxU
AMiMvBbKflp3mytPZYHRVVTWY1yYdO/KJlz2wQkqlRy/3df0LnM08ERKRh4l3Kpt
/DtgE6yXzzPGpe6svCOiO091YidmFawmsf33yww3644N0WCt2C1N7gLbSJpmL3LN
/RgNJl08ccYkIh0CVXsUZG3pOqjocR0VCA8lX+VMVLgtT1I2LuKRTOi0bqmdWtSy
ZGJpRCP0K5Nag0JNzv/r+KS40dQ8xwoKXqDYg8KiZp6tSRJ1BxegK8ibc7uBR/SO
vQinwh9KB7gl3lbZC8Zec6TCFkzJ9m3/qCwVCn8HdsBWVfsUDf+yBKZSCMga1ZUI
N/cXS5uU20NKPx0IlONRcagXaIyntQQu7iBFoOUR4LxXxW1PGNYcOaTJmxIWPNxk
CaSDYNR4xazliCOyCJ20x5lhhcLkOgJi9akWAzag3CCJ9pgUa2HLpHiOmbg3sjnp
d4bsDoLe+1LmgdQst3bDjBXo8DiVOW2EPmBPwmTEAPC0w+mRC7vf7OCOMipIu9w3
6MNsQFMtcJ706xpUuKlu1L+Hzkw8DESZe9iK14dmIWTSk3H7bNRxh7apQAXG4ckN
gjZvWPRIbtD8X+VTqKRJ4VYSjmvyxPl2n940RAzkfD+6XBlPo9dvSkuobUdvt8oW
9NjgmscjCKpt84Y//UKCad+SpU8t1+FZnITpOyMPC6m+uTVkcZBzDSYBbxKQXDxS
fccqgzqExH6flzqqnYuct7zHd+bujt/mVfkq89GShqFJj2OTFmHBSQp7D0I6CLQ5
nwI4JHikIZRC6R4H3VsjolESkU6MoQKZWmTSA0sQz/Jo3PQC5W8FBDdvPY7o14VE
kvGVHVem64Q9dp0AG9WmdSV52UKIRuwF5iP5Xt9b+S2u0EUTi/K3gYcVRGXmz6Ev
tW3gbFVea9pHTzQSYnbXL9bsbRLUXa+DkWbJM/ZHMVJ6eGI4uDF1/qNNOLPqiIYk
oGLuYqR/agz6Nx4ICjEn485VPT6xs0JNdQRya868CxQzWxRtSXak2IS0RiSGVEVU
vWM3gMm8qFBm7BvfIx39ln0EolmJECgEczRNgipEkfpBluPm1Ohx3k00UF4saBql
C6oeHzvk2l7KCt2gWuj3z48B/ZPUlDpAR7gzyP73kBSjC1cf2FlisN2uP1bL4Knt
Jtiw54v2uHWiv33TK0tIgnX/JAj8GkbYqEM4/p+rwVRa4Bq7sXW9EPuURt6t9yIP
D89V+9HJcPL3hhCKlvkDGgc6znQVF7uvJlg/lgJrgNSS+lF8Tf6zQbaNSo3FELon
ziuZwKtgvLNBBllZvqbSa59MjohffSE21u9OW0Fp4sszaKqBHbnZz0gwU+6Mh9Uw
KAtEf2mMjM82psGDL3RfndCTv5III2BTUOvWRDWuk7KKirUHKPoGf8dOq49o7PrF
s4D6vOALuv3MCNNwnd6FV5Vd/aCalgzhjowAtKDDAW12kr7e+m9pgYKur0NFNrH/
41ft79WtQlGGFeI01Wi1/PpwTXnr5VGJczQL6y8RKsad79LBZqbEL5JeU/EUr3lr
QQ+SeN9XKnKqxkp6iYBMtEtGI3T1DWQCrRz05mKJyyCd4qqp89iAiL5uoSouueqt
+w3dGODdXN07AKHfYQl0u2q8eBVtCdRPkoU0Ah8Xl0/n+vQSPpz8G+S2HOZze2uR
4drwyS6+DXx0PmcJwaliQKGaT+BM7GHxJG6PpSK4yntGTJ1bTR/FrjY1JGk91QoT
lKKO0YawdORqljaAYpt2CBwOKrGSpRzMWqqxS/EX6VQuOx/5viKRqbHa1Jjl/WvV
LDWF6PfyxmzD9S3CdLWIOn7CCQLVdPMS3z054xrOZLEzW1Qq7L2QJW9hg6UcAGUX
8s156J0IOLGBBzRZU7mkUhBXKZLGtfMAvcfsQTTkN72PxDhk/1fn/9V/QTrwFYOJ
kR8w7KXrdFngoNKFIC6S28IuZ/h3mtJMSRixFksge617Pl3YtNgrOcoGaVkftSiZ
WiEZXYpBJSuDjlJ4ShnAn9x12M1vPqPqTGCdaMIDjYO0+ujwmdVAx6Z69adO6ci5
IEH6TexbT8YlnDs5jMWtyEldzKLQLbIODSuBAqfbknZIyWJnDvGE2ZaKUFksSubG
YriwxRKJT3egzNZUVfjH7qbEwksymrIs6ojvtXloqgmK0CsD1TM3DgXUXpYbTraZ
tUsNHZfxuglhcmDiDFve+sgsaAtlOj7qBiGKcmG4qmwlXBTpARLYLcdFPRrTDXoC
m4nH0oHFojK6e4QlftRu+7Q+fwnFlclNX1Hil1Qm2iNY2ZCBVO8D+Pz6lg2E+te/
KiULl9hnJC2G3FfhwYjorCuDRF+MERnEeSohkGknj+bI9unexCNiLw45ODKphm4e
xNuG9sSzoYU1WkWwCNYWMPNrZJ6ZRVBmd52hrPrzQuWfWXY2gHx9RVNjRU/ERXMQ
pVRD58x+oggUa8VduXoBPfZhhFS+G0Llnl7e4k5MDAoXduCjzvAt++wrTVa16w1s
mwtHTvlBhTjNsQCXEw/cxTxNCiuDX2ekRiLgJi3ya1WcD/lQrLJMjLiy2DVoj237
/XjvszLfCKRy8VlhXkaWOg1jkEq01pVQ2nvP2+9JYYc9S3l7olDODqCi6QN8vCp+
6tTd1VP/pFagnd57s7mlrM124bDVW5YGB9xMiljeNpLVaXvGfOjApEFhyEh8yb/N
jdWA4eGgDalsgoc4EyWSwZVSd2dPqxol6hS74XToisnAsHeV7A2BIOx7SNbxC5A+
QWOgwuOv5iuaZS1He7iEoPJE2kmizbmV8DYMTeNxBrtHapZJLS+YnjN2vEcEQKGE
AZdZkwDUNjobEN9DkwW7dffW2LKS5tc0nflm9BO91QgBhTYloCAh2+lPu/FuQJFM
506+0Z92dYMRGdS8rjUCsf2fa5U1AKSOOqySd3VM60Qh/A6cjuqA+YmEf85YJHGn
yiCBaBe1fIatztpB5BF0FnHH23a98dRqo+gppzyDAJ9ATrqKuiXOWNXdeXbjqsBp
ITcCQFyU41vlu5kjz9knqAapyS06dLddnhoP7tCy8YGg/v2rq6R7psApiZW90y2J
sGWJobtIfa7iSL40IRvsecWKTBqP7b585N3vTFj5TVFm61RmD9z3wLMHHiRFe8IZ
sIuVK2O18oHEiti349AZZqV19xNMflVhMesglEY1OAYg+1LEVFsSjZjacqYweiNX
OnMwgdeav+cDhQLgGjHoe5m2AuoXH4ZrtFc1aZTF5FF7bxty1D/SDX9vl2J/izCN
tL855m4lU6JI8tNJ0WEcyBoh6CqRiTC882+1z8M0DGdmuc4cx67HCTM0NNx0W9vj
P2ZPWGdYzj0ZRHM+LRysBRea4qUy0ogzF8JqrryCnyQt2Ia4vCDOGyOQRcKP4Mfj
GO/E1s2PnAPYi5ToRmYivSSlLQQ31ixqNTzCZXtXmfqjGmPx+NfskTQ/FrhqudfI
KSaqdmnBmaxs+VrT26/g2gDNn7mQ5coxt5dKS6VpZHhTOUk2a0eG5PXRdu97UtUM
p/w44XfxEeS35lGQECgTgiomvY74MznIkziBZ2v477fEPhPP3Kskvjr89yXZcTmS
DM99DccuxfUtk0Jny9BiYysOzEn5hOCDf4t5vBexdhBbH9KWcyGY/N7qsHwiYO2J
4P0HI1c1PnJ0EcmqP5pibyb/QYi/OzfS932Q8SjzpCcs86VvlzaoCPSAhFSzlp0j
5UzfUUyIGSiLTLixlmDfIi0JCpRPu5D9xUomtUfhzPPCXEeKxZ+CWNBLJrSXJEtW
E16d4kFp5ASY+0YAAvC8mXUzsBg/+XyxTnzW0PsJNNoYOegMOyKM/NR9iRs5N0ib
g2WlHYKcFBb2yIiIm5n9wdlP1P/qLhXfhOCM5J2vYl+Jkn+iAN+r2f05uU/8vp/n
wu+70pVq/6Q35z3YWcy/MHoVbFMK4NDB+DL1oKb0ZK4zJ7Lm9BNKVLsU5X63bXTn
Mjq+qM8Bjyn+14k5HIBXvqzfDJGPvCLEW1ax0nMdeYCOmNEeuRsbq1N5538e1x4C
cbQu3UYtLX1kmarFKQYde9vAF2tzyg9B44mxNbFwFPbDXVDesxfW3SuD9SgYpVTE
tXHLsS/FMQtBJbOVToW/R+2wwQaF8O83lWv875cFuwS2p8xQY5FepwCOlZX8UMRT
y6iXdff6ecd4Cdh3v5NIvwSh/J+3dYt+Pqcm469XaoFRwZ+jX0K52tEaAR+g072m
HUkws82x1IN9Jqgf8OP1sdgsGbkp+ui1lzMlRuYAnwdS0UIfos5CHPR21hMFaeP1
j08Z2qLgQy8St51FFWTjubZ+D7XYj6naJf+BHB6KQR8yTwyOci8A03d68RTgNvBF
ub8SLhb7cAAvp9DS+rNzPZWYw72zm9gZwNXKaYNaAQsyn4/nglza9BHSaGX//8Np
ZjlrInG9kR5elHdhFRbyFQHA4rakpLK4jiy6VasiNuvaNJfp/p5PBv5iYJfyD1sB
A2ZHp6LIbyL3aBGLAS8YHSpqJhKfXNx5flkyekmbYLipfVh0zJB5GtmeCMkD7sRD
5SejcYoyyNe563tNU8tgUuQL3hflVYkRyTJSM8g3YggCNHIyiHMNVuSKMJeHBjIa
mzJuPSvGSU6bab2D9qLcY/UXfJjnqASdYvv0f6A3GoFO/SbSt0s7lhG17Tp94guz
eQ83HYFetizTpKBvUrOzvi5BZI51j0+tFg4UB6P/nIcJU7ug/RfXQLkRaLVmFIft
SQtdOGyEIDFs+NG4RXGsiRjq+0LRtIJRdwKTCaAnV8ODxNFXWhGkt2h5cRzHelBm
bvuXyA21VnCdR1ntFIWsEsSZb6ulL+Ff8DbqqmjejfA5/4OGDC3KtBHRQ7pqZ0hf
oAd7sGmrlGBurXA419yEE46z3luKUbaVturdO0Ir44jSHQ1ptDC1stiTPFRlr4XK
73OxIAVTUHgd7B8OE9Rc60m81YsqfPLyjepNDkFsPftd4oUlUqYjqbMFaRb178o5
GCcJ0Pl5xVBgPt62hh7/7aIsUkd5Rkdp4aGQn2sUT1iTwQO/E9y1eJJBW4tQemOl
08oPTKuX+6yt5/VclLce3w2YoCUZ6pgudSQCgTEnes4C8wq0+KuDGkUOiHBOjSOs
VxoT8xSiCo++ONJD4aZcNi1jdcG536sawsLLc4gjwBgfJ91KVWgrLhpX8od8AnPZ
nSzKTbLDG1WQ57Kwakm4qBOaB4UURcB45iMHCTuSnbfJ+Si1Ay6x9Jc22OzGJJYi
a9zmn9YVY+zTi45jPhNYmJZdbhg4QQaa6S0ehYTZr1HCXFNW4DtinP/mu1s/JLW3
8QAhLreSwjT2mTqRc+9iibhx7mFP7zNL9R6/QG/BWXVbOsT1pfjhvb/b6tf5zBWi
cl7hp0iJcadlQR5mQerysdExMQwt6xQDyMFo83pJgbDwgzwyfYVUCKnef7p1Zrlq
raeuX/Zv3jblVr+fzhEwdCwbaywEUY991NMoVyuEg9XivYjB+M5kniY7yY+PY+Nu
efw/D5N+Ep+xSKa+od2uLmWHNtnywj37x3egwDhkAn0/KwBI44dAy5QELubJsNa+
B8e5JG3EJoDnBxRW04/AlrIxrolb+cMSPnckJUp/t0z23+YBnXTiEHdA3jBGsyfr
4NkDo539bOmUhxNvithTiWxke0pvc96VJ8p96rNC7vecWnD6GujpPNWbStODvaLk
GjFY/OA5C+mEQw+/rquIox0j/ZS33beXTyH5mz1898hVvckbzlTnfy3Rnekv6U1p
39jlLnz0ZDJPNkncxcgF/EIp6R8CJ65PTf2gdGjYGq+RclAuc7+Sy5h1w4n9UDE1
R59TLqaBZ2cCWSzdwxLK0jPS2krHKsdhciPq/6sAbscPec6upRjZKBT0Q5MFJKfA
l9Pvp4VDWfXCEG0itqxhGO5MdJ6Jp9+KKmrH+MZqt6FQTa9QRtdx7ZVRc1NwXf5P
vxz2bfvySCDY+Kz3WxMK0/zUxepmROr8MOJDtid/l/1HjXteykl/PyCOOY3FpdpX
4ABIAqW6bC11X1aKWq5UAcSC6Ersj6856nBOKt2VWU0RH0RDugRNa7ovTgk8oWqh
0j1muxD238+o0j0aK4LkNMKu0okj9BVGmhqTgQxCkiHGe9kwBSEXlCAEnXZDHvGz
BdkFJo9Vdobmmo6teT68duFLn8mNwVvHBP8sSVXO9jXFBct1rbx7Spvi2kq44JTp
Y0kzWTts4PQq+RQxv3B/vG/po1C+v3deQS/WPRxTwxmfFoDSX01FGFjq30HWbKRQ
J6PsC9BZ7B11ih3xEaA8Tfz1V72aRd/gFysA9siXZfHidCwtIdtDSSzBPJfqSb8n
nK98eVJ8Dh76qyiHhUcstWV5ExfTwqkC1P5DSAVeCJi9W8EJS2QeSjLXSFgps3g1
nigcplubQQBhjL7uFV4hGP/W8DwhdgT4jlV3FyayBbEfAnroHDNDFf+CGUrs3tiJ
oY6e0lIVZrE5Oh+ysk2s06mKopDoydWhkPOfLrAVhWepKVg3nyvT+ZWEFHu/kNQS
eGsfjL4CUmQ0dXaNEh+wOi1Gm/FT0s5ci2u1stMGOXN4G70KXkNydp98jWO5dG+O
bRm7mvtJUjieJWkvS2lO99fq6qXSQMuaQU/5rB/5yXWcqdAhl3kYHkubfVyQkriB
4xndQAhXzUwGiQAUrNZNFv5mfr7FYRLNk0pDK8myap/MLVsu+9BLMDH+7u0Esdy4
du3Sc90iMRnmvKh4wdssMKX72v8yNFLVVogB166BR2tCzTIxOonw72Wko0Cs9A29
+v3j1Riq5bD6amjlj75uCt/211hEROFXgmSvAAcym6S0Tz+xBRU+zg1bUVjgQHgj
G7PkT4yv0Zc/ky8vq5AweI76LYer2hIlRGB8gi/hTirlZUxNHB7gBgFqIFmOA1XP
TgRlMDzmkR9GZqFIRxeLDzJGdB+2lDzWT8agV5gi7/zaxija0q6ODaaZC+QPsVpQ
ntAv9Y50EE5/WpG8pLTORotLkRLeQcwAgTr4UnT5jgffGzXKubRcPl2D3gLr2DxM
wmATZHCNuB/z9XqJngByoDJsgsJG3xl7khOt4/yDpmgucdCDfZZ0vFHlc+ruELUe
GCf24ON+/t2FWOBcdZI8dY4a7hhDiYtIboCk94L8jA0WOYyL13BuXo7c2p9tcH8v
WusAILdrL5vpMpFpAkJpd6AIjRJkjgJIgQpLK/PZKetfyuP2BuhqJI1V62SOgj9Q
O8WInEww6IZ7t/fbdDZFkoxHwjTrHmDXC63Wa1ANovWIVhtOhnraQz2lCh75prxc
soU1aHD4aS2kLdno8H2f7K0QjDUUDfBIBHoOwoLf9bPnJtK+Yz0418pQX7LbsxVh
e6C8HRqKR4M2JDD7EJT4XIdThue8f37oV9YNeJ5GFRThqBoGrd1bdLzY3GYAtR1f
XvkQMehDdTgK5zFdx0o3ZIDZtL9Q7LEqJR4GUqRaInL8Gl/iq3ZfCy7p0yw1f6y3
2BBQjKpI40tWCVXniUPqqy+pl7TNEhQRiVeqZl0oA8fl9wmMLl2exz/rMTCp5N/q
CzxrnUB2jkUFogWsN3EhDWLcaKGxH2E96iwnpa6yT9eaJAHebnnM2zAf5Caza+ip
Z4XO/gdqnfRMAZMvGHkWqUJUiTYGeF38j4AXBcZaI/AIqt/PPYhFhX40F78qnmlD
FPH9xouiBa2/lEYF/E2ge5d1YR8SZbEQaStfpzcZxGaiFOsI6kSPAJgQjKexnXvT
3j3wwhx6vEh0FuWA/3bBiQJAmANyM75I6spCiSNA8SWrpIr6s+bunBCG/nZZk4Ja
L1dADX8ywYYFfnZmPDw95kVQTcCnlED/UFNcV/Lc/nnyF2Td0PU5usUNhWRhdtJE
BFXIkewBqrJWlFeRPZ2J4DZVja+kYHsYF+vvuuA6wzuWj1HxIf+vAAzFdwP8j3pp
z21XA1rn+Css+3mzuQQ+/bJQcGMKvEPjmMJbWF8PPMpiK9th70zgXbvCB8q7Qtk0
arBGg6XNvU36ASwPV1Q/gv9B28J7kKyXQh5qyHE+waWZ1SCvZjnOWbyuSV+N5uHp
rrEfFr/NQ7P9T6lChVvs1oMZyG2t058eDmG5JllvzUQ8I+egjgO/08AoFnt5xbPY
ULh4s9q/EQ/myETVdujuwSU8sYQnfFAGFFya7jdjltsRgwej3utaoEGx9al1tt7M
3Kcv3csXIuNir79j3n7hSFbluUidGdYHkLFuT2S1sdUK4iWMplZ+DDr2LDnsm3RH
bz7HJtvNrBIsNkCo4jMTifT5ep64m8/ZwkFbpXpSiJ9n3bIPE7qrMCRvrjevEHxh
lR0efpQjd7a3dQyaLnscA517BmRf6vYvkB64GxWfIosezgCwaVYk0hqnsSjs2YwY
Ad4jQaZG5cp94+V+b3AW3nMQHWyi/C7ZAy9V3FgTKeTyqP0lHqI8ymn6112NkNv0
c6G1lTK79hrX9PLbTdoa1Ngcb8c6rGimXQvB6ooOSxgUDf58/C2pQgKrmZiijJN+
AlcPLOVJE1UQYwe+VfMCgyIilxrjSQ6j7STA0052oKISpDloBQTwixXqM71kaNyZ
9+9miKTJ6g0e9rF0taKHt+Ceq43Hgxfy9Yh8PwcbSOkkTOFEZcz6xEejpTNESc9i
Kp36AGkjAMdR5jLKb0jVKZB2PZi64FVPwG4EpwAkTSsdgLuhVg+UxJ5twIeGvQW+
sf6g7eeIY0WCojZa8zHSnPIjpXjgMy7VXNssWej0n5rABMDnqMilsEgG4LHVdTiq
8XHqbYzJqELlqdoia3n4Vd1fLS3hKKmZGkcxW//jQ/wZLLPouzJaKU1fiEe+xARi
M6M8pqkxS13p26aiumoBITXLM7k+mKY2fLuJA6TtFFkIoxAjCPpecvM2se0mH/rr
ST3KVxeMvLkgAiAY5cQAE7DGaJroJrNe9ol9o104yJtpZcbwVgjqbe+JLOmzpWwC
CauM5sfNpdcx4QnTZjNJPf7Uvg5UDx33lmbYYr0EIb5ccR7h2oFBPeVvIcMlN75R
awi/BGZNCPCkBy3Zs+kNrM799SHoVc9CzMajRkX8JWFzJV9lrAAKZM9PoJ9mFeI6
LX2Cdm+mmWkEqSRDz6Z6DClUeL3YA21kGZ95uODXAKzLtcxtN+Z3oJLiub2klp9b
yQHr8y/xoiiwHV+UChw7O9DKD+lnvYMdc4JbrpggGE7WkQostiA+BGjMZPfIVQcS
6jJz63JNY/JZ85xspv708qEzAKjtJahN3uzqjAmrLwhPtL8qK3w+qq15B3NF1WUM
kWHjiRvV5ZOTrIORE8dTXCVhC6+IuQNjHy/1Z36A+HK73YJjn3zf1a2n/3Jvbc2Q
r3fD8KPOBjHlwVTQ4MYWQbciPc1sHA7eX4p/zA+xVVo2XtvFNbYWRoO8UJiCD+0U
q8y8TAZA7wJkj9S0sDsTCBHwqwfnT+dH60LMnl73gk0lLbg44i2MSPCd+baBQN6M
uaBgYdB68lAzIHTU636lZoIrkmDYjqc31AimCFIBsrfhuLvgV8HlDX3paxlmy3jP
LSNs9FK65lGbcOIbh6hqKWxGjbel6UCeYIOD+dBeomYkd3bT3pjH49BjxiXCbF5N
7++XdY3fxRVGEerpzwBi4sbF3LlN6A+KakOP1yEpq+VJLAe4Z4nJlISrzUBE8Sjr
qZFbWgKNqDdHDJg5EmR1g50HD4WTeNtZVfmUjg+BS8qOBOfmXx6SJsksQtCVzJ69
3KLpdKEBBjsmpDlIcaI5RB/65BWinXLPd7K1luyN0nEqnc/+H9MQQEdvbsWIySB+
kZDA37818LehcSwuQatgodJTzcjlGYbDrLzXpx7HmQJG2ClfFUg/ZMvSW2wEosV3
YRehfN5WIb5njQgQS8d4Zg84lft2gb6fP97cWlLJ4+7QIVhchLFpaD2JdcumTbnr
nr3iVe1/jWgh6RxBn047CarvQg7Zl7KllacIDV5nek01MyqSsXLiq4ZqLBsnCkxd
YC843T7l4MFwJp5okH000quxIwZSk0jcIP6UeGG1Ok1h2JV8qokqAYgF7LFoFYOw
y/WroZ7eKfuxf73NhipcLX7LQ8+nXy59kXxwmr1LIYS2ruZKKPmCBJrIi5Ou2MMa
IFZKC/Opod1ixmJV8NLcLSpnqpxqX8Sf0+NekWAEuNT5Wyzzw4Au4kN/XCRCcO6i
ZNNg7OUHfjmvPW0heLd5XdNZ16nTah99BIvqJDKWQ+VVwfvd9gHoiagRfD9oRtnu
n3Lz/QpR3wDcZFMnf9YKq7BJwxo32g4HvEnzno0js8thHa96jbaY9Sakw49fVuik
cbQzyTTmliED+AUxCJJlNBDHX93iSwWzf17sMKCOHhOcg5SqGU9QDIlwqRQ+w7/T
kyAwEGl59mhvdAYsUJXI+UqOUjL50q1AeDfUgPI2a+xE1tag4DdEH/Bu7jDM+Bs2
0PBoSEEYkmQVGabtiyliSt43/hgRckcaDvUMPQybD/dGosqqKW52jlJkShhMUQa/
4vMbvupO0Q0RQNjjRT9DMPzD0rVnq0MaGarwtkOxlmix29d0lvWHg0vNZg0HpTcT
xuXy+EL7pNiFi+i6WoUBx6rJEtPbNsAW1nWAJcz0PX+8aVerc/5qQoy/KDGpXyX2
Xg4Q7GBQL2BAmu405b/TWyiV9hQlcxSzFQsqye5E60Mqai/8nkvmLq5Y+tAJJ/Gk
LJUmiM3lxYy8MlPpQ6J2w+B+CBUoOD8wyqB/g9yOgTeaj2lLBWHUWjvhF+EABL5S
CYQaM87A3Ioyq9wX5UFl5rGAmghynLWWoWVQRQ5Mlo1hDJMDdoZa0cehEOPro+AZ
u52Wixfax/AH58z158HzSleRo4s0sYDKLFpl3e0bLRFFUDH81QFzG8eJxrsBHkYj
qxsjcYuUtnxJY4n3IXZoCK0pN7OYHybwiA9MieT4BATmNXOh+SttMDL86RfcWojq
BOtvRu61IBlRpb0pHCtKDUGUR/IZIBEIusduGwivxO+TMw3j69ov6crBLPdmGFoM
loKCg6rK4az9S1Jjrs1z1BS9eHv4J2O5dVHMxp0DyO9NC5M8I8TA7JDuuTILD/Jq
1f4E8KmHtmhOxmJsYH9pOBXODadLGlLnEV2X5k/XH4NYxNBsuxXyZCIE0MxjlwpK
IxDL0weXBFOgJRTt1uM8S43OihKKbjPLjnBMfRVhOYnART7uSeyPABMgLak/6AtC
funF6dFfI4sb+Ou9YdTuSwna3+jXSje6Hh8t4nr2Uz9PnXC4ZiqLevGGVqlv9/QX
BANrSiAzdzXVaV9ZrHQoHH1RNOuYrzS83RpO8TIQ7ySU8KIJ4EDCZY6LIVbKy4/Z
MMiB/anEzXpywNqdBgoQO1Z6Y/590+235CzOfvSDWpsDdtE4IuPmjj+k/EDS1U8V
S1mA9lMDeEmbV55lfb+kNWcQ0Td33E89V3T+UlO3V2MyjUwavQqE3qgB79tufG0r
ap1uCLkdtS9zocjk7Pit46VqxUiHPj9z7Lh9fkFR23OUYjllEn6CikndC+QIWNbh
uep8mBiz+Q2hoLe23clt7FBMxkYxLFGKl9qoMm1AbOFw9d8FWozYyFth1alQxe8Z
7kktkTsYa/TFozL/ADWFdsBo4mcWfB3H3nDUgcuPCvzHxW3AgYxlhfswOUgyRs8+
epQjoLWJec14e4XbeGiktZYfs/sj0tbZlPDqZmdKm4Jd35dIsfy0pFzVZV4s8nvW
vTRVz1J8awRAAVn4M0WOdfz84P3GjXVFUHlwwjkUwF3UyWk/NKRw1pVkTBhnCfMl
QWQ6o/Er5jXTPum7PgQOJrbhdO9IYZ08wZU1vw2mVL2qxgrPqriNieWiIS1Ijty2
MdtUIusxMjvrB1DixaaVsnXgIu4B6WgT3mneKZO7QN8sthtBj9hgE5WdAE7/B60L
Y78Nk/9mSgvhsdUDgN92688nH3z5+BDLp0iQaur1HDeLduNN0mW79BWo0pku17Oa
xqQRtNEq4WQ5+BfHw/dHVtQg4SKH+4jvAFP/FUomyegbyWcWOJrCqBDlpMbvp5gg
zhiNYkhVilXDL35qrY8pjQ++P4R43PhaK9XtKIn8wwuadTpQIez9waOaxBzj/MJk
zfEn97h7+G++Zsr5zfXP/Roe/Ft0SxiBqI2/WxTq36xYam1M52gczy8uEG/Xtuwa
T2gQbO/wyHyXV3l6X3XMXLauQFuaeh2pgA6/nUozwnirnjnITEkUqruslO1KcClA
v3tdRrDYrFxJ/Op1XTVyWkKgn9w/ayAbyf0+yc3kb4RVBKm3AVqOiSgfZIUyxwbo
1XIcD2348rlragiNxXmx/wEYJk96jC/Cbq/xGDGkSe+scf6/6jhNF/G7GbFBgK4o
RyzIzkYK1VTpq3hvlrG2s/yPxKsgz8EmNMUGP/pJAAESbvmgD4lnP5+oW09PnM9w
wwWlQtCwDAnMtfQD4x814SPOlj0m6OwZg/FeEnT6jRny42w4NOIJ8wZvNAWYNQDr
j69B7C9Xny0g+qY9trdVdhAlFbpiSiDu7EAQdpjuVNW8jXyk3SJvJwRistq6bz4M
PeXU8lKHqmX9MLZMk4RymL2NLp+Iw2Ig9Y2JrYlrP33kfcVDSWwb2b/Wo/nfstrQ
iDdXropYb4oDTUzghjRHVsrN34LA/f8IL5wDT90d0da4Z3ZLx6yqwqpYu/3SKT44
4TDBoLDyzMUpuGRNE5gSzlPlIWydtQAmwfmlx8FPClyxpzz9PkDJQ6r1PUrZ4u8k
ajU8v6URtFpamclgU7snO3j8OVKpuG9Bf1BO0eTQTBiO7ItbqKjAPQTzQJg0Uuzq
rBvTEYf9OqBR2Vnpv3lNr0kiASg4hdT7W/Snu8MdQ9Ug5lWp55d91KCQDAdJRbtb
hS4dJBOMMRiRO5TxXghM6zpbvmPFdSbk6l8MaKLp+xpasVg9aromyLqGlOJGoCQt
sL972cjBVf62JcxeJLjsCa/Ol9pd5Jx+yeDvkDj2guhh7eE0LqZNvZpM3mMLEfn8
MdXXJDmCzVtNfPZtHMQwxyXzhTxyVzeDBtdTjbXMYIqCeeybYmIwM0XTHc3ibfzB
PkmAGa277I5d5AmxhBFhsNC8MZcEvCnXYM1J9bAt29IhXLq65kl9KFpsgH3+X/5I
nujOj8IoSKWldcK2p0SljrRGjEvD7gGZZLtG4Wx5+DDIQa5jnOA+j50fepBc9GLE
145stpPxHsy5NZNRtZijo++GbTYIUUr+RJB3KTSRe3C775XDutt/FvD59GQfsmyG
V1kctl/D17GZki/NvWVwOHmvfcdOB/FQFPwQVXuLikUi+1Ly7Pd9oEIiy3KOfR36
Pxn4Z7Keh5mZtaDdekQtb9yPrDv3CF42JP3/81gQ0OC3EQ+Q2QT2nFCUlb1yg18x
KzdGVwA/T/+IgR/wWZN/ZUjY/qKXsjLCgToRBKSN2I+/+4Cb5FSADtfosJm3K61Z
27GV6gr3OmnKzBqyKmX43DCdKTDJWRzmFIdQkwwwksnaRDIL8cqhxDawL4EWjvv1
wFx45QEiJS7qET2hiheYNV4S8auoepdkE1NC26102BmGFFgUl4GZZRygeSRX2fy3
APeLdkCBS/aX2KQp9fk6dmC2jMLWwOEcRrv/W9p+LwEBckF05+d2ZLppE5vDsLZt
NAH/rhOou+Ot7icwZI4FhObpGsST30ax0gp5HUSyPlGc44I4pPpRXNF7kM4Va1H/
cSM4niKdlhvNAuNatOAuCx0ThhOKJn2f2oKfnLE6jVLRPPjjjh8nkJZqC9KZE7EH
oypRYU070pd5/AK5fIqJd2tVUiP+ibh9F+ynJzznIX+Wv7ssi0NdE/zMTXnTsx1R
29jql/49P5JgpNk1x4j1wKtnY1Klqi8VgrLKm03cmFo8eqErefgNkPYo6+hWGiND
ATqkw6DYatU0jJ/TunpJFSgrrlGHqRMxdw2NKgLi+X+t4XoK+GaPYiC59xbLdaa/
d98hGGd8caMIwU6ZsDw13zsZhtDZ8CRZ9gADDDwkOGXQldK+EofCd4WgN44zrxZL
n74eVq8acRC/1WEyTg5TF3iWJvxC1Sb7TTBAxzTqOppwdkMSDvxytUAaBqpf+VUR
7/cD6zhkUq/5LprPze6JeVDcn26PjWtOwjFpDrn8e/Fdkh42DZC1ySzRUAEsBquu
KTKKlb1+v/1I1wK8weeIXuWawk+ZKqeuVXU9vT6p5+WkWE1Rw+Ax+KBG3wyDqXbO
VnSD1JDlDjrOoOM499os/HJ9+tLaSJ0w9eMY0zUYkCnwpdGOu60HYQJbCpEY/uQb
iaj12nyzaVWwkVH51sA5++IltLUOBCLwO5NEg5URpU1hn/vJaW3dzWrYv4fxT3/a
YaIvl4Ljxm4sTa73TocFU5/rcrm7CfipPgjr2kQherZmQmJweEI5NtUGkKKz9Nh0
SCC+rpT44iCrJukBWiaWV9vwfuhhqza8jgniWIX+hyeMvj9zb+rnvBElGX/6mteV
l14hgOP3DK/uoNBOnUrpR74+5sBgDwk5lpuaFqHh04NVslzuMQ8xAESoQAm6EJxI
Tp/if0LeJgDsjHRzlxvyy2/4fVrQP9fBNzBRw+O+b2LYbLQENWG4dfHPXOwpKbzV
tMmeBuP8SuLtjZCVKcNVNrcWNfqqPtqobvny4lNz2UtO3qDyNVPWO3PEMcuZxOTZ
QaRwdaPd7USU2nyQydjwzvb3vMo4gBHxl7gFgXu7zyzXT+8dEooBfTcYNextxTSk
9UYwwcbefwupyry05HsMryVFN6y0dM9DWfBGArBgXEkqwkdX4VSkLE2IiJ0vsNmc
4MfteHqJfoRwQ56gsHLb4l3FaCSD8Gb38iRyqwwM31mEisZfeKp/0H47wKW6wb1J
OKVs20/k2h3bw7ijEj5Cpz4yzjXI7W/pAa5rTEKQefytlCCdZg/mXzk6P7E0mzNv
eGYHI+IHYuDMJKn3aJuKcx1jZzWX+czS7TVAFS0V5A0CFuFQ3np1ng8VT9vSVakx
ctQE64QapwITUTGDD2fwis5VAef5R+YUffryAU86b91267jDAO/pNAUqv0W7IFKm
2BkUjsf/hdCOYmSHm61b4N3KocVI6Pdp1CVnUmRmsO2uTBtLO/pG3/T4gGQmug0K
nZOqhxQlFYCzMgX1BMAJppS3hUmi4hI+6zNBcaRmIZ+rNvyICN9rIoDN9TFtqT85
qs5UgK5CrLSiDa7orJ7lMimiIkQNLDmNbz2Ui6qrItAJphTeXCqadc9GAfE5UyUq
nJfHe7yzu58Tns8hPCiYGufyY77RNKJxmtdphtwcMfnloPK38wbyDD7I9YYtcSsv
1RRh07j3T5JdBgBF1TJjTQRdoMlhUawqdMtI8aOXGGmjXzG7CB1iXHxeaaNSoRfv
Vf4EDyZ5Xqao6dXms2EEfg2rAS+h0ZEYBwH0U9bwLiRJ//xTjz8udOOL5HvXQwq8
DHbI/B9syeOLRZ5EHhE1k9O23gGcnUxu/AxuUzyyGom5UQLDoTXxtxm/EmZp7yFN
fOAj/zDnYn4BGNccjkpixYCWg+iiR0+DZzYsMVQhTxoVgQ6MqkTMJ9IaNdhqJ0cb
ZbvMMmuQleO/EGVDL/WnvcyNJ1qJ6i5s8lH9Gxql0oLvbxnUySWLFqBN0s7YLySS
oqaMlWE1aqqizMKkMSJjAksrYI2HMQCM7yw1I7MITARl/7gZBX7TkgL25ekyip0t
/42LUbVbF37kB7kQP80PNi7J1vGAsuIzBqE+7FiBy0+cK9g2f/Ko/6l2L6amVHuT
xW/cmSoAQ0R26vXESU0RXddzf3VWDac/hLxqdpYhMJ+BVHQHusIU98qcoq8lgxq3
Mh74pbXRurDCmCAkLJeVm8sywG1ivZ9pFaw0GSOP/6dakqUkGlWLmGoGjmgHdPEi
mHTEvma7mmIG8X6BQiYTLb555RZoUHMVm+Aqbl4KO9piiy1E+JKnPQLDZ+Ad4vRG
GP/wINB0NeeOKPA0Uho/hQJ606+Mrm3EyP2R8AaYxmg1l3H3knCAfOt9QipwdXbt
b20Gx4LsvkTMXhmbU3WOk+ykRn8T7v3mwZzfYYjRzzDyUUtEBDmTvmyAON/embzt
4G2zYsxrPp/FVAIPV86fAbS/S822mveH+us75B0bh5oG+Upq3DtPMQcFeFw3aVpT
6//vv24T0L7zkm5rC5k+t2z4Th7GEQtpGUnAS7hnUCVZj6/5e6dcbHBBsSv5iksw
nWALBNY3FWWpYE1d7LimLCuszfH2hW4w4RRk4Fa3fOThAS7xW9z/s+DQNvIubK6J
W3MOFOv7oy4SgyZy4Fil1DzgNR/YCR8Z4pRFvGKF57pUy9Q4Z492/8N2bLzPSoUB
ukuAuXjtHUe4f5m7F7UxPSB1Kr8+HvwqaWS5iucfflpXywRQk+YuMCMIG6pX41nB
EDP1mvkrPTYC5r9oeoTcN3zDhzkyYGp0jIB0FjUofbB72aSc9liWqsFPJfPDLUhw
2KeR7DwomfjtQyBZYt9YWPs7Q3RG7cTRrZqc6Cqqg1MgNo92/U6r4LhGYLFh+bh4
5GuxKS+w+6W8ux1lak1jR6dJLMH/e7PgBshJ/y0RizJAl2iGcmWpV1AKsr08x0rx
AF14hqQW255c002aTh3YowcTUc3jwSmN7T0WOKuYyqjeLaE+9MmZ01eDlLZrhzFm
OdRBT913SXVdG9wIGM5GfgvlGzBTARHM2Slc6X7SODWc1hw2t8x75iBA/IXlCRhM
Z9A8xHSgEk5R2JOePJ2PUTjTepQ5ZCDqeF/SaKwet9hOKJZ++ltQ/0jvJ0RDJnkr
0tRjuuvgHX8orS990MGoQ6PUavUymu00YCIT5QBT1yFjo7q5OSRC0chgcpD3wtNB
TeAFwb9JxuMPUbAHio9o8duD4tNVwsBkG9k9AW+VA4kPzz1iDZDysnVABf8eNo7Q
CHnBcm19jABxd6PYOx2PBHBo1vZuZl1VXLs//4PEOsSl/7K8QVwHZSANPliM9JSq
EUFB9CCRC8BhpSbPJDN280ytr6zeOb7Lw3oCnHS/GX2+Gfm2ASzN3yOh6EAsSOYv
WZFcqFlDczGd/wQHuJDXidasgx3aSGM3CqhijJIMtLqRnINv6Nhyh7AVFru2aX1t
teSnkis1Gqbrc0Ppjv1EmwqE505/YCHU6gAYwSxksn4mg/rVrksZ2zrVZSe2it/z
AYGkUq+yk3vej26IeHywiiVT0V34wJz8U+dFlel2XD38ufOb//N+XeMTVeAT4Lx2
jXoxtVz8Jyq/Z0N9b1EkkWJ//908tB91/MXm20qYHQ3penQSbiGRwqkpLOs/eEq3
Xh14p2IZ/IFie7NVrxDerbGhoGoAn7ZQwvn2zOzMnv/q/mATMMuNsLVBVkimQpwN
aNhZDGZATRQ9XR/SvhVxtprideHsTo4gNwrvFnG01lUcni2U3F5q+BOxAB57XHFn
hA/+9tIm+wWWLzNHRjFM7r15PdSf3bKNoCH/OY99xyHN+7Cl4N2wUyAtv58Tq/k2
Ze05zxTwL0650mJs1kyFdF/AlfDBCSaJBh82fsYtjYGX33qvFKw5qW8+Nq14j8V6
T2QHdpGem8NJHgrN6Y5S1wMD4xrqjSw7Kw6LfWUX3d/1c0oLkeZdgxKiiBylMLxh
U0HkdwM6L2mjjjEBJKOiGWbJ5Ur9ovoFChnDD+k747JH3diZzqzTh8nrChQzXndI
nko1iym8oAGKLUbamSo7ElcrZpwANPCu2AWyiUwLaR6PA9GuQd+9fyZKuwYs8TFB
iT7m56B1DFbiXdGcp6ICMq6VTSjEXG2435QYvZb1wYcQSpSGYY+c3+Ym7fo7mzqM
38IdPNREn2gGo/sMGfgpHTk+jlTTor75sdntowDXBTtAsgoe6araCnqNwWJ6+rwa
OoMCmCjOLtAsXkjou6JYLoiwHkmMVCCfrmnfkkZ6zSf/8lztydNRCpgA3fkceM25
+P7e3s3jbD/gK0eWthZcPNSf64PeGVSV5Bi4SDEBl9TFQO89NNUOUUNFRRS1KJuM
VyfXQ7A70xfBlzFuQWuueq6huEPAIU6dvx/8q91kVr+/x6dK4uvDWV3dm9PSXASE
oW5AWnVIpZLsJxnnD7B/GaJqEymMMDkHGvzlRp97aXLGSu0D7/THF6smCxOCDdeC
xK12Ofyj3NfLwfv8i2HWZAbuZiidZ6TyqLeGC74HFsN1+II9/PaGXzyGOVOvyNBZ
gwtELujldlbst4ybGRItlAJ74r7ydHBuGNl/q1FMD+o2KqmgHzMiwXMatUCvVCnU
595ILANw0PPq1GCFA8UuPjzucIFLgjqQtplqhoJs453LdAKs0wpNb9hR17SRZF+7
a+PGTAuCC0BaoY6ShVOl+3dSnpEiKbWpXu/VRkobEfMyj6HOcUtJw/NvRWK5/mUR
MEmeH1yynf0psRqZniEdH0HUiCF8CUxNu5BgDv/Sv+y2xlLQn/EwZ49CzpbT+zU+
6Ez6QANL3wgw/3Xw7qdGgVQxFuQe8fXziH3dCC1lf3goSmEABh8O3v60m8Rdk5Uj
HcSUvPNWHUJ4yAABpItUNI065dCcFRG6hK1b68IvEV5Da1qENEF5+uYLF5HsNYKm
JtecSTcZn1I0Uv0uDnrvxSZn6jEr6EUZqrhpVi/1fg6tLtBXUtDWl1GTCEPwXalj
8Cm5y35ISkDpu8k1dz1GR7nQ9f7DCXMT3CaPMhbkyBtPjaVUWekqf6fA4f+Cisoo
48A2RO5lQyoiBqJMlouDVUAh5Z82MB17Pw/0FOca+n312ut6bCmkcXcl7PB0Avd9
1iPRow6Q0fVeIkMMhcmb/YUNFCsm38c1wEdTGIsgo3h96jeqUW8MnoiY9YdTBBUC
JxFjwAP7Gz+8mkY3OJbrFq9y7cE4Mr9gv10ofR0pEXmjQ6seSFn3ZAl8gSezG+XT
FkEnvkqshOkoaUw6Rl3gTNhAF355fCTFLf9t+0m/Kbd2nkLi9iQA0Zd6qfL5ak5X
7DpmEjHHtk1p+nKg/5m/FOM3eyjhxRW2pj+LAGFfe5pbAGfPHktzE+FWHvLMNl/N
3qNA3vgXjJ3wfKFyFMn4973jYCwLDRdxvVzw78SdrhnWOHg5W8sNG2lX7WG0KXWc
W+xjtM42J6XlrO+o0s4qhcv3//Q/YOlBLJ3aW8GqJ6xGWcPF2/bw2Vbe49MMPUUx
7BeGIBL2zcUc7FrrjFiGnyQEq3z32uB5Zw+T76galz5eAgweKM601jKqsfyNLItC
Dtm2OueML1hQXXTQEDjzn31bLmZ2OJd1rXu0u6m7LqvuFH4feygo3UmzcywDgXPW
ZdGeY3SMzOukbBOYT4XAOGACBMz4vU445GVT/GX5RVeuHyErBgC7QkFj4+GGZHJ4
Gk95ePVLGTb1xVdzHCe5wzFmmwzXToxm7Vm+PAKbn9NDty4473m4wmY8iworsyg7
v5AlQ3UvcYWwbyniL4QegzV/u6IHt5RlYZ9hEsPuC7+SwXJxQ21YNZ3gCTaZdvKs
a3eMzWNUOvN1TxKDAde7ty982lBg74LecASNIS5eetdYOHmWrJxr/qcaodp0rJvs
BqGuBVtByQsLfQTYdxShbBcDB9wPwsSUSxxBI2F1OXhTUO5WSIER8f4NhTbpYBpF
39VVM5X1ARakdu1LWhNLJKNjA9KNLM4s9QqpogtBZAawW1zIZbTcbt9bTJ0frEYr
g3EOU6e+iMtcWYW1tY25y15KejQAK29HkPlhkExaJ87TjLBn6eNdCZrG8sestiv6
wO30y+km57DbLHvtNmHehGjxCaMH8M+S/ogcWmjtRLIkXJenvhmsXIuELSNHk9MT
35OMqo5g3anl6xsDN1B+lHtfI3SKgtn6UaJFmclr+BiBfF5t/VhmLVvTNTk8Vkph
BIDEghi1CnclypEeLYruboYw95Qf+iIJH4RVT8b4X1jhzhOo2J8Y0jJoJ/Pzhu/H
GXnfFgMtKhvl7yXTbuUG8syfd4F+C3xTe9t4RPUJkwf3eISXivvOrujxDu+ISMEw
rCENOyKaozDkiDiq22v4B8NNEjrZZUJ11/ryDa4fXpLzjU/C88UN+5pE8RP8hMU1
QTKppiDzwrCP4buoJM0yIZ9jIVypNwWOB2ngY5yNNwW8kvxDADGUu/6kxCRKrSh+
BmiYyVhAkasBx/LXdBtzxPP67QOE9KHORsgtShuPN1zR01ysuOoByMTvToJythHY
llUJtuMjIDggbQ3/h9XTGWob5gSNz+k1uTv/WSuNIyoCI/y32cP1JNIXYyOJj9pK
/mMSU8lx1dYiOREQNBd3ECw9bNIe0Bl3rCCPbzzt1HE4Rl/Qyr4RX5zQYIkKMYNt
XNOG+qZ+kIvy7Y64+vdHY8hnsQbGLuslS2fhAUEnYOnH+WHtDvyL/OF1pWxd2o68
0mIIMs9JzxlBhgn3D+qLQk1DXgiAmdJs9igBaT4DwygBsb1MpYNx6D7ZK37S0wMe
9N81IA6fKbOt7Mr+AAGEsYKPJz6YgQ32kgK7ciD+cpLmg7xPr/y7HCXCykUZrvob
35e9zEH9hgyNiBX/jjDWsXAI+lL43wFAupvNlVDObZaA0x0VF8JsQlyp8L/h0nfO
RL1a5kxKu6Q51NLtyCeot9Yvl1ItQiEPm+XZYnQU1vNz8ZXZZlQ5Aebr/N30rulu
7v9NDk3DZIxnUTiKwy6/NcpW498PlzCRgHYjVURwJ5mhzCUPSe+kg0vXaaqPObMI
41acHs0HFiUzctltPjQhsyJc/m+VRZNt3i6nG2dNG3A4oDQqhscntaGktWEO2alr
l2wL4OJiUs/Eb6w9G42ORPHtE9N0SczaCtWXOykh8is+/wWrnChUOlWbkkCqQ3wu
iVc0zfUo01i/cbf269kVPX+fHuHBH5CS7Ap+UPTtOXAoBwFWC69eUMawrLjkMygt
EbexDUT97LOvuYAOweG2GiuBf6Pq5yka+7YFOXPVbQgc3pPqaWO9gqqm0q436JBW
yaGTaodLRKQ5l7ZCxPRfr514BM/vB4cPowkfd3DXwqM1R+KtracIAYDRJCi4uAnr
/YnvqNZVKSzHQO34+DLOepTZ+RgILs1U6Pgxl6SMqtJoteSq2BofVmY+X29Q2xch
xwQKkW9pJqdA+K3OJGDubyCWg8mpDEILXzjpa8miYV7/yq0+qra06n+VgNotS6Y0
/PIwehHb2ZyaiTYBlmM1Pfr828oqFeQiHU0+ss1wDQU6Q/BKaDUVB9NSPb5cFqjK
mOmyPJ0I8SDga+JTH8miIsPbd+ksSU4BkpX7Xwp7oAXvJ5T0PDqJzjSIVWc/X2UU
31ke80X/TDIWk5+JgjGKrf6FeNC9ZIsQz7JkMgcyGaxEw9sjlMQIEUas7/Fx+caE
jQu+OAuWzrJiOufILKP/0wayaLjAu2Ad9RTWb4iEWEpbO54fyWDlCfnCAnqoQKDF
j9haqSIaCSjdQjdLmMg7Keuai00hULieihCKHgRG0gwSxfAbbedbQVAeXtCLp42X
xPj+asHTgUeZKPFs07SlW5st29dsxfoKnjmQ3fA+vJ2DeThacJlXEgtWB19Yv/z1
XpGgbHaAbAAuGhRRzkU2trb6T67yW1sZNF9Mi4qe79NoaQuDp4nT9lFM9uXpbezQ
xTBwOx1jkaMF+lNmzUqJ9Oc2vb5kV+cFgvTwbVozy/DQaoaSVUj9p6n4Hy17MaiY
9EOf3qEDWXEp8p/iQA0UJEFIBtC6ZvwfQrJw8hZC61jZHDp1C01hzRFS1JDEazNG
csecEVtPwg1WVv7ilt0SOENDBM93W8UFpon86nao1bGBoyJehpkciL37S4bpitrW
fylL79Byn6dMGCxfP8C1lx/ZisuMl08QhEJwFBgerTz3lpdmuAJvpF/NsXQvY/oy
W7jPh06PGqFW+Z5uDmkCFfeqp/8t/r23oDnqe8My+QdSn8A41cHGNGjrDzsH0nvi
J1rGaDs+/MxdPIHF6WJLcmKytFHYayO/xUKtBh8B2aH7F5RNeN2azbErRaQSByQ/
oMbkFBDBFEUx0mwgfKy4Wu4g3XXv7Hk6e/GjLhlowYUDCxUficWRz9OweF+JNVfk
nEELJOFEnZiAbaE/cEX8VsgEVQGmqWSi5MOErA78M722mIqcIYyj2vgZxyhFnz7V
ZzH27aknbFMXPnTKiuUD5ahEQ2pETzT3AWhBB3q9GYZ5Jyjqznk2KMYPGrwttBut
FtgOU9eDrXWSa8gxOD2QoI162dFxTa0gjpIuuui2mawfNI8HtG3Xds6vgTSaCMyt
6WOxxyrBIi5eLcRRjXJD1BxejErVqS0G/7mSdqbQbPUVM34HwIgIdCdPopBuPcea
hkJ7tmy+TKiIlI8+8kQ4uXgI7o2Ziu62ti4lqYDuoUHBIv6vlaLw9WAI8iEbaqYb
HCLFuQuIwFlVtQcGGUyg+pJXY/B6QXqousjbVhBYyj3PB8Mg9OJ4hS50jaOdJVoS
XLVxDGjtOAj6w9L9jI/UXnDMqoc3NZ/PpBtJ8gBroea75eahqtjcloNVBiVngRzD
4DLSgHWDxKSRplUaYfYiswW5P+3O6FBB6MFkGmBbfJeyo4WJ+TicLtWD4s0QwQ6T
nF8kKWlajLwU2jSQIfq/3QJCkDJ50mvN+yU8BwaBYaaBN90nMRZhSHXRpZYZDG6q
O0hQ1pRE0qyxJkKn05WmVaz5o0ZxhR6J/MVckH5onuHKXVpZ1m8AAqxjh4GM6QuD
2pce1R5lNxsU0i+0fMc9NZwf0TbEA+civixlW2e0K7xLqArsEtkB20PxMOk6kmYl
AYPNTFWwLUa2b+ItsXxZaUoUHcehSMlFgxjyCFAl/Eu7U8s53OogbO6nAMfpKD0k
0SOrpDv+T0U798kE9wC5N+ET/K8Z5I0JK8VjcZ26XQWXT9BsMGoZtaMvHQ/Rr7eu
8SIt/L87QXWdABvUe9xj0kUZd60SVSsc4ph2hESp21ZDGpb2wDWw+Wm2znrl8TQ1
Z50Q505BqEGnefb6MHDCcMWwslmT1EiWwg8lr9rxfYRLSR/NMRkZXQnRN8iKs2tk
raqXcZJQKuVSya8O63a3WWISHv579bsdFzgk3U9EchZkLRILDhbPjNjFq9p9yzgL
WiaIqt0PDZ0eUZ4D7Fi5tT1E1qR3vugTOGKx+e6pQqPOLIb9srMGOU3nOpKzQenR
qh6TwaG6u8pcujEEOdUAlFA3rI7hSx91ZTye0DMhdEGa34tzsKf0ux+/jfE8lcWl
NgvIp2ZiGmael6IxuZ/oMV0SWsl22BDD0SUKCOvGZfmQ8yXVAVL9cpU/yPSw3GHh
Jj3TW7THJH15EdAqZ6JbtxiweOa+6mrZrRy3uRwTQxbDZJP7c89k6AIPqBZeTJgT
Fm3K43Z/cS2z0atFdADEBbEvHJGzvO33eDBFxUnGTs3kqlnlBK8uJfFZSRhlAQX8
6lIvMcX+bX9WEb6hkEpsT2DffIvHUBTzh+vkHyMwl//oJaMjXZ41PbIxkVnkgD6/
SRXn4hdTB5qWWxxBaQ2RjMM9X4EkvgSUxjI8x9SGmIUnGj06Ep/sPI4XNmenh2Ky
+rWDPi3ERgrJp3Z97TNkUk1rI3/eZvYQ8FoO/X7b16p+ACLrRd/+GpWZGB4D4u98
rtnfGWbKYK96UG6Yo151tfACNewoFe3ZWtklfAcE609wdrWYprbFHN13I/hUZ7is
+sdbXHOUJIHKUU5MS3V+KPV8Me52VXEcL60JzSFu/Yd5IPvCsVZheU4U1dbeqJZc
6dgPgGVwyO4oTdcypBNqTYSc42uvrHftCCTDcjbMhLFjUevBzqVFdj5WJB7nnWfk
lG30Xa/YRt+TUu0kR35t1wjdEgamtJQV+a6QyC9Ty2/IXfAwalr27mE4CUWoiyy8
7LiJRgRbGh6d8h0s3GqOfvO3kO5ATEDn1ww82zKTUUHrf4o9sPynz9Zlqlr3mvSV
+O0CFdGuECpDXYqncNgN62LbSKvWUhL1o9ecWyO9a0asEN9t50XMLmoQhhPW6kWT
2T32DYDxfvqiptYN2YNgt2VifB+yDlJ2YLbB0n8aiSvt0eKHIuZGvMgwhq5LGpHb
e7oHI0HUhbtw5dKG1jthNl9zXj7anvSHcjHpG++hPhJGiMpEQtxNjuImVySSlddQ
KUQ+FzcIoVFkciISwW++KQYREpLDWjLX8ZEvwdOB17pcUFQ0pbEmMeG5bdc6H0ar
Pj8M9jpRNQfCu/5u3GhRGa7gHw21XW6h9gLEMpzOrEOkrZ+tw74OpW1yUKAIuOJJ
Imt+wiZqxM/IiYXUqQ1KRg4su8+jOkfU5K+qM1hX7/GfvUBHYwWOFZsI7ShDRmbY
apZeK5P2DKkNfVVhBaji5zc5nbq4+by5QwrziQrwmFh8pXLGKGKCKxEiP6j2pbIw
ftJ+uFCQzSfMWPa0nM5NoOxhz0IExIz/ZdvdYRiZjdFPsXT9OisAHJKnd9SPtcJv
fzxOnmCoQbPx2xkJZ0dHm1vSHXpdg+1fYr044Gf8Q6PTnk1UPvCZYfRMEOSjAHkI
66K3ky46vHVcRz2S252ur1kbq2bB1Bse7dTgMmFMv45cJ7afhT+2c6g0J3onPvSy
41iA/4PAZe5b/LsQX6fHBP2zByiLsY9b7pNNyw92hs737oCIFu2Y5At7q28K4Rhn
NRzFozlz2q6x0V8fD/nrcpxBmNeRE5GUyd4U3r9ED0P3aDL7mkb17Ug8hXrMLnuD
h9uvql04ASVRinm+Sq8dn589dpK6TTZHyhkoRxIH3S1x5PNfCc2uobOk0zXlxs4Q
3NNcwfJ8OayT84piza9RAAKyiQwE3ScjmVT/6es5tcKWo6fQ3J+cpP2jTBM/5OJK
1udL/rd/WB1B7sRCYiEpwe6diNX/w2qEAVqWiy5lXMQA5C5FyQnDfdNzCIsdpw2a
MFtHa6jRdkNS76BKlDWSCPV4y67qgZl16CE31gZaxHKNVAZ8MkLK9Tv275NwLpV0
z/2FQIFRC4KgdW+97Wr6FG84h8NvGlUt9ztjOgJm6NFw4qSNp4r5Mx+l/LM7KbUN
W1VSeT91V0aTSZaWJBIlGy9Aei94bwrNotFyuGw89sHJqihd2V7zNTWivE2rn+9z
8lVAdCSHA7Z31AZo8ieYEo6yb2qagu0fvc5zT/+pRzgTEf/cl2gePX9rq2y8UEzr
M+CsgIOpD9um6WkE44vpNPgV9CnTUxT85JvGuoDoKEiYi0kjKPGi6Hx7kw4IGYHQ
esdZpV9XFhnNS/DwlTG0TpPHfXEITJnwFtNFRMpbXQnaMG5s/PipG+zAin6S6lXs
6BR3ovAKI9RwHKF5h45olAS8QQhXAMNpMQLTyFatRTuKKINfBzGRa8bQQRmYhNY2
K2d6r/Q6lOCvUM7FKdxp+A0q/NR5oRuVKs+LQCP6ZBHfFjyQeTaYxo1/ZpY2VCKk
7sEBHfv0jMn0cniyh4nvIQ6Th8WW4+rPdRHT/XyOdWbeOu85DxR9JDOBEibHFdiP
g9B5P1aF2P8+ACEGfYL6tu8DFC54cr5EgoU4WoI/FEQ6sLmH9xwgq/kAdGL3lORh
+nBFFMaurKhMceLW9CfaJY3w6v2NJDUt3cQDjywRF5ptXK/j07aB2/4Aow7AQ4Td
P7sBVDu2btswUgRBTaMqglVr9HPU+Tt4PbInavYvOBdxMqHNkvLnXKl5FaitQMGn
IJZJQfpyQ40YOGb/NlZUpuPiylVEX9q4o9KOj1WYPFTZUvddD4HqfXITDK5dLVFD
h8n1BowiodaMcOCmdSOzkJ4eIBA3ZNc3kY6Gi8Y8H73f3WqyKjRu9tiFTOVIfiMD
mmUbDyWzxtWKGtkV3q0XbxpzKftWstFB9PvZxpA6lNo6KgbXzTz7Q1xH+Wbhc0uS
FhG9CHeWSajFpS8GgpeIbMnux8hYFceWRzoL9n5QnmqwwVh7W3B6FsfYil4GgjtJ
KDowGZ5LA5Ne1Ly8liCxADgs13flXLzGu2XC3nTgBtHmltJnmWJXgyuD2Cdan2pX
KsKD/e2d6Ja8X9rkTyobD/kcz1DknZkDJ/MnvkC4k33Esa7lrNR5IrQ4LKrSrAJf
05Cyulq/ISq4LYGG9LJoZCVIUct2TWaF1VHncAE3po+AomDtTr2+3AlxbwgdKyoY
QJmwX940YelKldJqPhYBVBNayd3D2qX4/a0LvxCT0uBpftxbCp4XAxCMTCunwvWm
2be7k/CXjKFCHe9Owjwy+vVHMTlt+1HJb4AkjE6zth6VH+NEj6EYGKtnjvgzqDi5
Mm8s1O0dkv/40H0h52t6zRTZ2YNRV4h5aDZkXcd4r9s25V6o/FXTw23W2jt6COvw
vIzXcEyc/CtJmxu0OvUOD+zEPCptXfeduy5EJPccx1HZjvgoU2CAB0EtohT9TgDj
Gf4BZoe6frww/hUUFLFCD1KVM7Z1efzdhwxLoeQbo0kG+2IKQ/kIYrV+/Nr1fuu+
GqqWq0pl/48RI65w7sswxXD6OhxxapiN5lmguQ7hJMzp6Yt+VmiKwSAMW4+2KZx1
JpaxGzvAsukOI/yzmZp99vFYipsgvbGsmfqdl8a9ve1U0YVGpS24v2Y2wGWOJHF9
X6W5yceHBHwy4qq3Nywz1ulAQ1OW0uVBTk8EM+s/W6FA2ora56UxKXdOK8Xb8PHC
bq5qApfTLeds96Rx0T2yeW/DEhmrbDG+UpbqQ5FZbtMuFnk/5EbX8NBGKie/87DV
U+8GpmwY4tphvKYr1IrstnQBsFWakcXqRp8B7FY2qoqlwjD/aFKcan/gRzRjO6rN
P9x4dDRaJMtHBMTBPfFF5Vk+AX4TcusY2ZLn6JfnN3ooMGnGHo8bQX5QorrA42xe
cQYmM4bgPo7/thmT7KlG/4sb7n4JDOhXvnENx0htm+ncB95eW8mstQvVdbpRHFsF
Re4rceqewaz32htCr+G8gLBB3ilGAB0W3/XBSmCqM5zS1fWEYIt41kS/ZKt04zFc
ieeBHOsGIGa9GxdlqDREvccbWwe7Nk6RFHQQ2iY8vVZgYHRyPsbPr9qghChltFVH
fjI/tTV6EDlPrDk6UYujyGKDx6DadizXqZY3ugKa8WuYP0kFQnMt4CT2I8GnO6kx
GrPT7oLDmm8cqOCgHxaUlQ96leA43DYs50j6u303xTURbrbhAOSOSgnKmCe3/C3s
tJO20syEsyrDZ9t/xGGOsduB0+NzuEFpwxmwNOhdmin6oQ70hKV5x6dyMoy55tqG
XQ3QNCQw4Eo3Gs7m6s6CB1S9xRjWnd+L6m8A/UQWd05GRFqvwF5D5qN66RpTWql8
X1M228wgPDn6LRxSdIGu+lr+zO+fgxDLWEv/dOfPgadyNT4XYa1iyQhVq6xUGSmH
C/wlcBCAZOec69Qf7QtFrdGmkstaQW2HU5t3RnNQFdk7dh5xMhyduB7k8INvApul
0E0uiYzU55sRB/Q+tLE+D+2UnDUVKY4AVdP8ZWnisCsnXgHMCAmICvTiG2fogkTT
y6exDmQuWLIZVZcxeeaKSZZ6HUW7FkgZHjt422r59P4IXuFi6h1uWg7yv6BPA7v5
fLgNWLsfBhyZKLBUtaFbRn2P1egu8GyvMT2ed9LS7BBgZczBEvGUoJboVWCrpZak
n5sMhzQv3vRuD54B2/7JMwYQPWaukqWDwvMeJPjPlEZvX3kcDIxgS/ShArZMVym7
xrO5DNhOzenDiPv6BPuNYzSkcy26Xp0jxXh9ESK7GOnUfP6yzwt1r1tD2pK6O7jQ
4hGZieKjoX0cuD02IQFdQsmnoiarVeXXs7aVgyHcUX1PYoT5Zb78WU4Q9IpIKQoB
59ych9qOab2loKxd4ga5mZB3THjxN8pxdrwq1PibzB/eL9/mPVlDg1WGWhorTsej
EtLzWbjrSBYptpEKcjUM6UxLitvv2fqNtSpRMpl0oo3cSzRCSUKNG/eSTKoflFak
OOt9SY2xQuvflcLwLD8S++vTfOJJLz5jKdOhljHi1Qa4tG6qMsjcMtq689ygBgyf
H8fxy8xZi7Sqco4SXWoeom6lpjNr1XWVyQmRrJu0OXJAwfqTy4TanJe1YJNU0LpS
we1+I6Ux96ZDZ+vAq7pNmaG+W9trGQWh83GbrcYtQgiugfTxpL4/MEr6CPPXWhOP
MLEGiED75jgdq/gMkEj52U/yu8cUbY+9amD1yUAkNA2ANxSiVxCzwXhCzW09Lvu4
7fDnWYk31F9HBptlMyE37YUonarpuuf2Ey3rCMn8XOPr3r6b2aPnU/fHlm+7DQxH
B+7KSFpWiOHyMxbKkdqaACYMSXY0w01XSymN55Im3gaCPx9lwaQWdkaFrYgUvRi3
uWxQ+fv+4BtfNFTt5+EjTVbtXNH2+H1WVmkJNM/Ly0pE4fsP0yR/YXUThO7/q4+p
6tMj0EjKR3c+1g5kuIaYD6w/iC+YZevwwGawbvSLFQiEzmpdHY6B+IU7srFe/xSX
cHVC17glWGfRXmzBncOxnV3aZ+PIVH3A2GSCZ99JlvIE6VWPlrrkRKqzr8QGsEsr
kDtXScDL1KxedU4TeOFMrXebkHpCVhyOXRZQimhZx5XjdrFDy88TDVgRamYDl0BA
4CPVi0Km7IqxWoi1XpiJdB+GWQ59VyHI8Bn0Rjufj90el1CrvrFlO4PjwddyBeQS
w/tbBfMBCsN/IKo3Kx5ddfrF8KpyXRThK+PLJbAYZjN2aoTH5XIu7o2askyzOW8H
Z39a+ZsOdzCCt9RrzWkHWJ7d48ORuhmKSHwwT/vVfr8RFeY0P1vIL3xrWm2ozqp8
dsL6FqwjP4mammj98n6hj9T9sTTefkNMsk5PRxXoWwytzrOoCB5HYEL2ckvHZRcj
exl1tdvEczMDtQGV6XBZHViTFKDEW4g0HnES0PSnVsMibtPik5yWengc+hqH3Qoc
W5fxfmRKCGLVTjMURz7FyBphy6dOJk5nLn5aYo7FvpcCKE0zHXwcsMWP/Xczf7FU
8nB6a6q7vWBEBTRU0kVGSGsFQzhXgmhnXICOGv7qchKuCmR8qAmXGcskuj2XCCJJ
FphEd5LEevl56KMj+zaB3KgaoPGW5Zd82/ohMKOyZHClzKMxiEro4I8yYb7fudT1
J64Pnyh81mRmxUih9PfjiTlxuTkIehoKeoRmtmjd+P/7S3j00hhcL4f4lOv/yD31
E1486aD5rQJn/l8q8BlL4ECZltlDhCQu5993AhTR4CU9/zbk4hNiGS/vUdMtb5Mw
M0DE9aPnYOLnoPvd42luBdye2ygzubahpwfGMTtumf6nTyKKrOC+0+/Z40hZEGMY
3krjxgjGkc00fyL8vQAqXWT6oibW3udDA/KLavYqz8uuVajtJ2K1l7Ju0uq0oyp2
SRO92aKDxm1oJJ3V5TcB6wxjZxbM0va4sSd6psVAUyFXWQHLx4In8Jy+LB7FxUBi
Rnuz8GbvnKxn+Iwi7fcJzZ/F9fWW2kLJvMZXFIE3rVZzFZzcWDk5stg4XrIh4Snd
JonVhhrQcNEPzo45GJlepU2Sd32qrHtdAqc24oqvRHIiiU/Jsi2jyIX5eyJyNjoe
VU+73WtwFGialfSypyRnUwikLtx9a4U0RA5SZOeANCKS+l+5d8fzL/XciasPdKtl
741kdUkYLitgjekigbCIRx4lQq5T/X3NPnrFAK1M6JBgVnD/GvW9RYvvoPmv+k8O
LMnrXPTIzJah6o07cfw5nH1GQjzzY8ZI8OWNss3NIxJJTi3mJ7GEMS13bZRJY//p
NDlDz+fjvxwaQsoovj2GL3T6mpz7s4A8UU5TpUPwUuR3G8+uiirCs4oqgAO6lDB/
oUIWxe1AJnPQLsy/F5w6doU7nCDDXsp2U8H2uwG27T8HJ9RFxJYE1SEM1XDEyz+2
Aq8zGcgiPpF+BJsIJbGa4P3fh+fm7cPdoSZLLEwGts8GY5hxyKIQUs7ix+QPAysC
`pragma protect end_protected
