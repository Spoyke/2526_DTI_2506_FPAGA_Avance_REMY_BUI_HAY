// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZPuZEwRJFOpmFw/abfTFB51OALdJtgKMP7/RIt94XDibTh1PGQqODPVaRjvyXy4Lc0QWqB3SF6JN
sjcxvH51lpyj64xKKhb5oS1YD9JaNrv0giqo93XhuMYNVEFiwiNHwz+9PrHbt8N1A4BqEqSBBp7L
QubSnAkHwkjWuKvdBSiYh707KESqREuLzHCjBO7F5XlSyGgl5glpZM+RA4lk6o8SYEMo3um/9dv2
fRp7rGQSyqH4ohlgBywBPUOIysL6ytIu5TgvQt8goeAubXQIt5P3iFuteyKyTACVUy5SNfYyuAN3
ojKveaIzQ383M6hXl81T7HdxbViga+m4MEeFkw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22752)
QRYsAgSxi87xWxPF34b4QHq0vNVGL/zN8klYCuoX/hGUdjeEMIHqRPpC8NMaTtnMvPpWZnF1rOmq
sPvcUBS8+k0j/PcOadpaKrwuXsCE1ZkIEwfKV/XEzbrRq4drcp8+574PXfb3V2nYBP6X3d0l6maP
CUaVcMZKKvVsKipYmbGIixcSFY4+rqtgsKKuiSQ57Q15Yok5LZtv0WDH91GCMALXsZZHsqwYnCk6
T9CqD0KSO11qLpNCCK9pJncnMzS2VCk6IR/LRDxpUPiSHddHmTe4S8ERJ2eCBmxjbB4yIGwQUXCw
EBb2TTSluIoJvV/sspyOUJ/KcVXcfTkSIK3Fz+7TsMPSeUeeZyXHmRnHSmTVUz90I2CV3ifQKFsh
UmHlOJ9rzPT4S5Y/ssGeQQ8Z6h13MfSf4vy+mJFgdqRbcAxcvKVIocktzyOR190I8uUnTbMK0lpZ
zBGkEHvQtUQhMYsuIrj//mUtW3F517QywAntbQG0MkWCwrkzUq9rHby2u0zykIryA2j8xqko84U9
O+AlpeDp8xF2SLv6q/PCe82mIrb8uvgqg7aryCjbffzyDDyjczdAtfTAbABlOgKrQzhiXAjzHZlL
8vncJf1BCMa3Qca0/oPw++biz8o46j0sIQILHlh7Ax2yw1qg0eXS2BRkAHl8Ow7XRGagXLlIlQW+
sk3RsQ7TzavLfQXrJl/hLfVPPUjKmFYWuaMv0Zbi9skuhiMLa1HudhyNCljt4Us0YfwOv5VSVH6c
6lK23GVXWsJQ8DOOrj4QT+kmQjQmOz5dFYvl0c9u3NiG3Y3pf6pkWAG4I49GCBit3hWf/Y+WssHC
h4YJIR3+ccp3tHJEt/gF3PWOHkpfbTAY2fnVqfas/H6znAWiLTFLhZuPgNTDgfMqqi/Pma6UX8vB
/DftfwP7eJ9gHdMjrXPDbwjrBrigxkRnBPtwSGfXoLTfnwD8Il2lUb9iG12ansRnFSkEmgUya4QD
sULdl1xKI6NuXRGCHdXS+UoSNf8Db8zJdLI6zm5fiGcL7en3qE4JGt6621EMP0gmnnMURKenSet9
0wSTTj/vtJI4umDjH9tEwU2/wXx8aCxpVvJBlQ0wiLaBPg//hzFZxIQ6BCnnnQRaPi3RtJgaSKlN
HBhRXSEyYTxLWdDi7jFTYj6qEmKRCKREgUpm0iC6a17rLgafr52fngW2JLVmL66wVVwfeEbuafB+
SopJSYUliNbG910+woS4hMjCohSFSN6jciVPizmEiVTp3P2fuHOLMB8BLoxovOjXzDGYzdpLW3Kk
xX59Y7OjfB25fO2C0E+hgVcZU3GtyTKvsJwA7g51+qKdOwB0elbN32tJUWa52GS8YZKG60CSItl/
qkg/UIjl13SPatkmzlbYx4HSr8P3+bmZviwdb5hAoZmgsDSQLNzhUysw/5xgM5dEmYhUMiZexkYp
StoVTBL57kd5Mt8WlYkGntrDc2S1HTcTY1jn1WOuqdfaCmFjdhZEVsEJHiW5X90efHljRo4TXJ0r
LS3MWBpT6A5cu0TWNeW5MXjmchax2P6udc7pgipGt+c6cbgdWNJojn/4qdm+34m/MxvtxCJNY1Dp
PilmQa2ur+Xfd+blNkRgSj+u6g6T6yg5nIMeghQWDmPwga2EoAVkwn1XGCYfNSjD9hJjjZwMxkpW
6iToiSJAUpHj1Uu4KXCu+O69r4BQe67m850GnXY9E0CkCYCU4vtrwENRceedgBO/3n2tNDfR3DyS
TlZH8akCkoHKoPb/Yka04zRsHWPYvtOr+HRaOuhFvyf+ho7dGIBdhXPBJPRpnei0BB2C4WeWD0Sj
dOKabNMdrgkHaQ1T7MQWyKxZsYsZaoSCO4D+E+gVEJU1box8BH0fws/KgZ5npAlim8og+6izwFwJ
cJc28O1vLFxI4WUx9QMSbIIKd0HWy9/0TfAJH0iX54xjjrDWk6roz2goktGfxwjWqmtZeQpFkPzB
OIF325YiGFZOpoVN3LOdAhyxzeDPihPR1DBCSaa3yYr150BHqxVsCiv5Y4c5XMm9JjjApV4NDgtp
THiLr/xkD9FKmZ2cNj0MNYbtk4ueYxlLyg/n+sr+Ja6BjN9kdp7DUz9hDfqdOJfw9EBHBOUhsiHL
hocNgS69ZS88Wl2V1xp6RKVOLDI1zRkeb4oToB67qZWPzrrWikM85yQdd96wKKw3f0QQVXrKcRI0
K/CjH2HofgbkIMqq4ce/H4yz1j1uvUc14XvxSh+CRvKmMbGrQ3m25pLnYdzRBquHSX9svJQfd5cB
Ad3/dJBtW7s8CLVacfli9BamQBf6KCLzNhTiNynm2RepR7GE0LmRkNP6Rvb9XOeZM6YgIT0YA4XU
ZZXPFAZMgxSuTMxzAXvO4NPMROjgo24IZDdWwX++LSiTLc0+mvZ90ZEsr4DxyzVAVoe00bxjmfWr
aYvn+xDWnPGA1wI4Kb4Q5RrmfgNgTx9fBwTRpQbg21XPlzqiUarOYHiJxoyUppqPtFFUcwyvd22+
80j0n38nGmTU4qqdM9dqLhtePTcA8TbPTo5N5MwjN+Fp2rOtxw3mcWtQo7uNjoE9yeJLPJP+Rh6t
tRHQW4fBTrbolRsMO0uEjLH31EQZozQE4M+ONHYI7qlF+wPIYSOrQqpgLjqhs9PJwDI/NJEKVU90
72et1S4Lx+9A1EIJ+HV31op966aUYM6LzzYs6SCaXVXKxiZs1GmMrzxs5rSOGAmaYH9uKacsKJKA
tD+2ZGOJD5b6JCp9x7O+pinWwPVxvbEfmq9JBpdDfn+xXv7sLxf61lKVC8VMVOFCsE/A521+peP9
Ni0IFM5zl4VXfYnB+wgGrF5bHuSefzCGuX1DV/eGdhOLwcBl0laD2d/cqAYKqqFh4PLlW6eWwEL6
0WyuPg2ex17A1J2BddF4qSyKzR1796z8/a4RTQVOwAiNtwxJeGcaIvrmKnMCLNvcYqKz/X4PiBcL
2E762rGuJ7k+dhceEnYxQfO9IS+0c2/mS2W75fPZovwRWwgZ0PKexHX968rC3/vhvbSxd17FJpWs
2nadTsjRXuJ2AWvp4/WSBtuHsb99NQ45Cs/mDrx72OQIkIBE/i9zv5tlmDglsFPHho91TbXmOKgi
ClaEEHAynefmHRgd+lw0mc4eagZLOCjUJjjUfa2HCoPhI666ogyTvCl2MTeBdtYxrkZPN9NShjcm
+h5r588LY0pWxHBQ+DfMVrnxPk6DtE14Y3kz9lBs6EFE3xlP3Ieq9JfxTQ7/n7rNK3F1WLTd46xH
jYR0IaZ6yiRYxhB1G0NKYHDyeRH5vclhJu4R+04ZweM+z4u/ocEieITwv/eC7Ri+s4PGg7dgIyoQ
RloXnx6wskbuqjoAiU2ZMuthsDbVfyf9NiMvOHGAPgJ7OBgTnPIla898AhINO3T+sFRxyVTcqgUd
dXlWNXkT4Kgpgb4vphVPdTsIPMHRQEujePkeR8YMBeGbLPF3Afb9xavgh6nrEtatq4elbtOBNlG3
sHa2+lqqxgUv0oGMptxwgUfass2RwhwfRbCvweu684WXnbd7R6mpT7VoEQ29L1CG5OMuJhWf73Bn
pil/IAoVAoz3kX7kkLM3l1m0K8Vh/1N60rj/3As600Q32dOT0X2HaiFTptYWOmy4R+zZ801xfZ2T
ozVzeAnlG/a0sKgY78Un39cVOFGOcawFiRHHi18j6gh4DEtQTCyL2BfKCVLT2GwmPJJrGMppw5nx
4K05w4jKLdZKOfO5MWgniRx30DOduAW3q3ZjrbBcT9J0Sy2bqkJZksEoBG7AksXnC5ZKro+2wdDj
4xseZRKVySJcKudD6RnwlRY2VezPYztf+xfz3VjXWSXKjysfzUZJo97Po+ii/ls+Pz0gfN9r32Uf
9knWf3CPfO0F6a9oRUyo1HxqlGzrmmfixaSDKbZXhmnPnQVax7FSyJ1HefVqgwRC2TZ9uVNrkGUg
pIGeQI391onJ3nYVcrb/4gZbVmh3/dX/wdIZjbB+fhrSzJHBWZnBOW5IZZa+ZfWDSott8sAYLnl9
YHpJvowTxH6NY/gr+OF9PoadMUKLldqUcAwfv6ylqNt2+VTlyOpQ1+gAFJfKPpUnzo+GEzJzIZVk
NZg5KUtAwmaPkuGn8ZDv5yb3ArSssCquj3RyZEbS+1uFdAgMjI63mydrpSGvRf/RrXsnX52pII/y
VwHpGLkFUWi84HbpqscjxngvRPAw7JP11XIo3mLxjqdahVhFnPW2R+BWr4kZokvN4Ybvors/Y0TV
uSePpBVu++CYd90gAtKjGPNSe4KX6lrzjU0SjOROGCNMP0RIV9IqYCrp8JUbrrc1quiYQNUK786O
7rvtEsQ8gE/so44qWs3lLM6w2YEo/pwHBNRrTiPhtdcKe89k3iBuZhTsn8uZf2KXpoHRomnqpYq9
upO6n1tuyJ6rgLqqyZQRDOjnBZSjDHpHIXK/wBiyfjw0KA5eP0U3xyinAZVHKeHEY1sLtH8hmmkK
tKcs+mG17a54q98UIMsJs3w4hz+5mBR5Gl3x02a0wch+l3KCLhlPvs3WIqF5sPwKYuatwVoHogz0
iDywP658uIV2OfAUfrQOyxivQU2+13+kQ26VNEOOBNjup6ochVocZK+JkXGS4RG/GvCmXNtuhj8i
5Fkmaj5uhnm/DhRlmPpZasyQgQCRN/fQ23aOjfIC8iJqV5YArl0XzMI2sPBnvoTXqlgNfAki9hQA
BDQsuC/yxCHHA7tI4hsWfrWgmVyxqcnNNRuqcQsEkPf4s3q4ATicgxdq95Wu0OaPZ9Urd0uDJCtI
wJ4VGLFx5tQdmk7yCWgDl9iaqIkxF9sFDgvEb8WfBN0tvpuoKhzfIttYLZTgMqGKoxtlfmE0CtR0
nI9erRCalt+DYeP002DoGrdZ5kR8QfypQzNlxqD6YcSbEmQCoEY+WcT1BvQ9T/xduxdRa8Ly637h
qvG1Fi/fSk9DpQ47NoqeF1UO1YL1JmsD1VjGqqmS9/RPn/VbQ+66KL/UdSF+gxGO2v3dxh6Seb9E
5PNrzjz/rpxTuns/RmFMF/8oGLlB9FKWekvWKLZeIX1SCk0tvW6+IlM/Ny9jj9/wImu0E636H2m1
0A/qZkhv8ElrLZ6o2Zj+TnDlOlUgIxvwHdZZh7K0f+3aRacpw4v9Jhh4OlAVw4xnayqi5SfIDaIH
pcb+73INMSyWRHoNc3C9HIEDQxOJO+ZatrCSLPROIL/o/R2z8MsHjjdAWdevYeWj2zS45Vm34s2z
x9jLvCAJORq4+su+c9BOpvb9XHfYOqz9SPJsEqmmLeMyEn7Tsl6mkekVQb8ZVnWHNawPz6Fi7DTx
DtFVRD3FODlmiPOVBRDlSY8mCJ+eHrbTlK6us+/nvi6rM8trxtaF4g+8krMCWXhteFY0Mw0d/Wxd
1WriHqozXskC9TgxQpTxp9JW6OGp0j6+yD4GoJ4tNcbtmgU9s2mZr2XIwDlHkm05u6Y3TP0gTkKW
cWhauNPi9OaZckHkGhhx9xeh/ka++d7bXo4XV8XzrIjaExQdBrJHckUWuF2iBYmAHhccGeaxcDCO
4Ijq6X1GbQKGyCUBabCm1/Ikyruc480fvEQcGe84ePDZ8XfSzd11LodkXSO7aubA/rRqQtYf05IF
w5XzGhJrTKT36D9gSfj4Ubwzoocg0GDFevafIbEq7Vsatb5Z7jGnKnhXP95jPfVc+kMHS/rEECRJ
E0Zx0hzZ5+rKJREm0LxmekI6mJZ/c77GHVa1kvDZwLyxfCvPs2dKzjfp6hxUpJtM0Q4eBq6MRCvb
Ln7avirJmEExz6tbYtdi7ZYxS+V08iDafHzop2NoXLQoYMSGem7roYloMeescEvmV4p3bd1pPuYB
gBDMlqCbB6LyutDUenoEVd2lJ6EQci5rC49GXhJygHxhlLXcm4WjYmv7lphrZikquN1S+M8A5ocB
Jpmc1dAq7fx48Lst8EHn7CbqcK9z5G3ia2IvRpgoWoKRTgqs5uU63P8EpAjIcrBNwVRrg+6D3te6
fXBcres1v6flNgCIWDV5ZsGoyMgQuLgI4wElJJgJr3qA/oWac9bOOFZVZqK6XSyhXCZ2F30YcJV5
jwaUp8wz40x/N524K18da8tHfHbBYdlENApD++vJbG4GYeICJyP8mb7ayTS//tWgbQI54f0pCzv8
B1PrwFIcyf+BLSQjjKjkJZYR6Bz0T09Ni7eVj9jMwZireKSqY6f6rimSDZbx6/nVrMDlxGkr+Rw4
GHo2nFlDoEV6qGAAaIcs7hqntzgc0wFjHN3kgY2dM3qlaNgJwkPBXTPMDLbJHgmwat64JXFb33QN
t5waenF9rJ+b/m27VYgDNy4u/biVGxojywE/R5tLJ0XFmPutoY3xhZADDHXkYi3gA8TpSIjBlMRp
Q/Y/6Kq5R/sRmWICvrh04YnnIItsi1EJf21KZ9auBnBnoeCbql7UzvJ6tdLwy9ik5hxRf4B5cq41
A0sQmLTHKJhDgTuY3KWeFvNoCvSOy4Zt8+KUiiY4s0NvcA6WKJsW7H9c4X9JbJmLQL99BTd4O2/I
owCBdkK8gZzpOAPcWoIEUshTH+E3MSK/KgoNF2udUbMZGvY4PryhsXU4BYSKydBF7RTBl8ev+eg/
+2DH4Z+VHqnNC91G7KArcpBsKr8OXtj22s7lWG6hIkYktM+OgfHjTOqNdA1+N7u+p05VRLlqs3Q3
ZPBd/T73L23Pld8sd36CK61uwvBEOXjTqzynmHp2nVhC9o3nyg3pw/h2Ib6DISnrMyy2BNEJ1PNN
VPxtAXZ3eoHssEb4oK7+JR/OELKRKHQR+9kVDh8XCWHt1/j3BmkLNHInbo/myTNd4nJiW6HXcqG9
uXoro0+y9mL9HF+Zh1YbQkaOCnH+3kA54eBFxHbmyvNcmpjzPwuo/Azs7PltQ1AJx8PVFztlXw+l
ROakbf7TocZZLsV1SO6uqZIomJKkedku3O0Z3cMivpY8T4KJq+hGf/6J1D7KVi3VxWakJ8eU3T43
Z9mewMPzIoANAXPXNx+uN8qknNX1N43p1BIVPMb59J//QAgtISd+iwsyXVlPRTiTXLliAQUJEDuM
AnkHDGO58ccaRQmzX3glkxNYQGTMGeKjslUTEJSoqWSIQzX6cf4YEgbblJBDBQSiqR3XVsPMF1T1
i0x+7L0IDvgyinpcLT8oKM/A3QZ9sec7h29AqMrj341WDHeOK50CQKD8sgaDGy5fkChgjb+Eghws
V/kdNwfcUbIcu2mA5Sj4UOwvjxzKo+vJkFLeBoFuXAG7Ck18QjAP+bq8v0n56MDy4Hhr0fE49zjV
3QhaW+W0uMC/54ivU9JhyVpKSVKouUwABbQT0RzaryiZx2UngCts9orkAdourRmOwwz2pg2SQ+V9
Mr5h5h1Efa+MkoVvN++Hd+CZ7WwxNzq1fSz3XDbAb1sqRKPINM/pwOqbsECJu0uRa83DChzyjPH7
uponoors7HJCU3MzN827K3tNqMdNgOSgHOX368uEpdUS9bm26Vw5EYwdmO6W5VyR2l9pMbdCXULP
bzGELiKX+3afnP+m9mzvewdIM6BX2ybpgctUTYHfIaGtMOepbryFHECI+SokHfehKDK7L2CFb19W
P+Se6yCy5xFM4dVZDt0FJ7c4ANjAksb9rumiKYykkfOqk8Tj0n4xdqYrnxcnqYF3vuc0GGsNz8Fc
nOLawnVDOeDSD2waFwf2CZGd/OTdv7D5/tr6PquW+foGo8qx/I2m7G5pGZmNZfiW6mM/Ypunm+SV
h8Zo18ilzItIoTHmAG3PT+yfZwvKwAbNBSHYhMXPhOu3yIenEoYspxZ31ztWoC5I8F3zWlPZXxHR
9YryU/iK8eZF++Qdc+6KLfUp+LqH2BFHrv5nvPCnNhdPX247G9RUgfPH6S/swvWCWyhu/zskgB/4
fIF08uCyark0IziktVXPHmrnWFJr0Rp0fWZ6+vf3j2r7IKBlyj2BBitehg6uqQMDak+TCXwROmf/
AO3FaWmnms80ISc5uaJ8oMXLmZcX7HLGSXTiIAy01jWeuaSkt6Ux3DP8m1h2ltpEPyELy8Mu9Sfa
9EhFtWmZXyX7IVGYZa654fvSeTgFMBLe/kTov9ZQqQ9F+r3NpmzTNax/oc9uhQiJ7B7ruGYGuZ4m
fQ71txcJEO4hdQoIAiyNw6mH0ToEGQqkzciu69f5mgNMG/ch20Rz1NM2y1Nr4qN13W7xfQ87rWPe
wmWFUWUGU7SB0nVhpsSFl/SJmhzeobTUlTs8r9pCnEiUhcJyNqvIZvLwMkNqKPeSXPIefED8GXmY
KDpt69hXidjD26fakmvWfvDbVg0ixeNgv6gbkDrvBvz5d9vv9qtQgKGdT51RIxQJAweNU58soKHF
4cRNniC3SFV4xehn+XE5Q8pXCs1CMtnmLST+AQxQ0/3aU3tsAvqyRS3v6U0rBF2WKfHFE6PbGP8F
aRTl/DYXEcrA1nj3rwLE8pcvw5iHHKpWKtjfVS1kV0K/TYiYJepUbzDj19Dcl7GrM4MulAtd4zaO
XOmh/qv+KMoP7czRchxKNMHEjb8XXq3bZguycnKKm8MksLyeEDhtwz0ZIo06xHPnL0WGm94eVF30
0bz5/Je9fz+tF2PdphLfsQLUlh2xQmuqHdKLKe/N9llONhzZqLU7ezl+QvFCDukqftR/hut/VoZF
HMzQvWChRIOgZNlqE1/tATfR4hWrNysEMnWAukZHpY8UreJbL91HpaEhLiIeSt3cqcfHuzUUbBrE
qVG1AVr7E4g/DS5iSIgLyFq49uf2dZB3ddNLNFieI6oazk0j3Zp3fHp+pGvx9H+EEZfXEzKmVj2q
19KImkdb+hFd0kFN1f/a6B0o068N6jdfypu9cnDXX2OaP1n0v67NiUC0D8l3EvoiDpwAgjaoJc6M
8tNs6BIdWIzZ9DJ8FKg3SUMmRl1fDfx/Yi+uPUfFZTca9jqqSyXUXJEXi2YJo9YOBKVw927MlbpY
YMrhrxCice0/acSW0v5OAcn+vjn0eTvuVMc0z+KfaqpHQ4E+8Z4UOn/hp2+qzLPaAlDneVNqAFy9
iTCiZ+SyM5ExySgjvPHHvYBTjRJF4KfPswxISLQytH5AK+KVeABtefoBXrBbHenxJAFZoHnMsaaz
iNXidQkSMTmh8IIarSSks5722+etsFAzzVoRXsbAUfYAIHocqcw8pAeO852zL14IbYqMnuKQ+ZJ+
GAPdMcrPvHDZtTMgRunkTEprgQ4jS2RFVrSlWQFvzrSzanVUExu/pUh0wubVzvQ2gL9CXnpYserq
rJbqL1HPk8aMcJ9Isd8NkRPmZTaicIJkatCeR65YzRP5DDl/HAJttAWcHPLgM3hXVvWSQICClsuN
/mLYyl4vAQNzhTusCcZYuf5R1PkJGoBnJjSQzceaa4Ndu+S+h4uL1gsh7t3kxN5m7DzcL85jm1Pe
o88Tq8XmuaThYfF8H18PuCLU/qIwhehgEB2eDr54vHq/wp+5BN6MIsKIfv1G55Exac7nY7N+70sZ
KvQsGYoSdkPsAFQ8iSzGC1HYnrtJaSNnfnd8AS9bPKSuSJsSkH94ejgDPp2u+kP5y1GKpTO2nZJy
rYoq/V7JRBmGuou5QxqAblDxYVdsYhb81/11D7bWs5gFViAXw4XOxhliDzPEq+v7pxLQ4xqpuqm7
J52JI6xd1s1eokEMuDWqNAyEGOgEdqk55KDN6BjjubcYUR0tAPrWBypne0mhQT2rzd3PkNpUmDd/
PIG1I2mAyCa6vZI+4xzNMkVWwxAjZDBDJyoqNNkEMY2xb8RBWdmL2rwC76JNdE1GamHmEhe6RkO7
eKvPKIXI/DK2AqiO7W26q/rfZujFFAYXf7jEtj5OWndPdvsFyhStfFv3OwTghBguTXZcinZ4E7Vy
wBpigjp53ak1qarWVZp+WM0jrJfXu6YZtHM9oRHIrioiNXwTv3NPE+cHf0nnOc53WBFSf1ZZNQot
a2bQbIARM2lC9w+EK0Qb0B1uQOZ009Ou4kRCPAtxMgqgaJ/3EaRUR7YQ2faF+9UjmBfJsKlckIF1
5wXH6Qw/hik6lfpzIH3eyTdwSBzYNCqDy1hjLiWZUyNOhZ/6ZR8g35+F68ighDXU9ev7ZdQollpE
vVxC8Igy4pgg3g/oX13AG/F7dHCBgpA/pIlbk+OhC3zRtjrnaSHqiTInBWutdLi63CchttsY/Yte
IhWLjMbXvwvTF5b1CUPh50wp8xuJD7pilw8PFOSibuT4r0ENb9rnK0D2Z7KyepQSrlxI6xUB15lC
/pIExMMYoX0niprcIe4mXScoSShBM/9rWanWtYR1EIANWFRUPGLRh0nkDJBdg+zwCImoiCUeTo/5
fZTQDb6pQhzmTarCXJQVwsISjyZIlIxYL3/WjATR36b1hOFOs6m7dn7wGv0OQ4aS3NW+klkNyXW4
gn5mGu0v+1oAZgzyGVJZ4LNVhzd6tHCoeczSXQWS9L0xJ9l+NJxbGpHrfarb36OC0uox7xKUwnyZ
zEfXLzslr45oM8vpjDw4/kgIVxkiLKh5KxCb6P5tIHWtbSS1PU5nPcIEWgqu7fNIXwbp7qoIP2D4
J6JovERpXKMdY2JJYcbsCKleLPn61XulCyrSAIGc6FHk85u20Q3pW4CfwIPKzXMPOFa1LnuU/el4
2RCTNRH7vEZXudA4QOwVDYR0d3QDux2sel9Ty/hZ0hNDrxMUa+aCHmBXienhfx1LPStQK2WZUwPX
JHKuRsPwaMPkmB85PZWFigeT4QvJYZ+nH9ctnmkDDmj55r2b1EgPGOX3jqrRtQl0aM4wfZomU4Ea
jPgRX5J4m7smkpBLNgIAjauPH/1L0MtIKmmtrfPreHjSf3YWOkEHKfE1BQp8mg6TCBpLnzfp+T5V
rrOdZwev3a7VH6DSZBsDSv+FB1TOHMYvFE8nMHoihdAUe3y4z1fLj4Hsq3hTnZBGWY00ckNvC58F
/jbSoYDSNFyxFsQbacREoZMt4KqiIn7wPAzz3UQLv75lSer2vd6Yir18aN7UATMNT+ZnVpNR/enI
Hovmu3BN9W2MPQgiFuj4VqWwo0GaKJ/H/lMnZQdi77CbVOAYcEET+QUaop9+bu6CdjWyatdeZ4OD
kMiEpKnY1tD7M/cDNr/e1N//nCqRlJl/8r4QFtoVLSghiI6reGmwXCG6nq1T/HlxCKp96RTDYpXt
sPzvHiPpFcPZ3t1QvoVxbffbZ3Scot9tkO3HTvXFOP2gY3A8jeSOOjPU6mTyNiqkwdlRT6QTg9NM
Cs0JmYNehn0nJxJJxBef+C2MRyUIkkriwsCLGjUTarCmRT4T303kXnZd5t0nt8wslu+BPs5fOH6g
BkFp2Gg+WsEODCPohRk0cPHWOp94Lkzad1ZDX5G52Aupw0+5I6jTI4W4tQaj9RisVAyMQ2Rfjgr0
bCHLg9Nv2oSED05ZpXspcq4c113LvCz885x7NFqqMkyJTOZKE9mu2+hnfjF9eSm4r4K8N9OPulDq
rLTC3X4G+qMHejiuOgW5s/trFU9LPB+sUP0iKo7TwRsqW0e+9aV4RMK7GVQgNnJ0mu1FoXXMFWmO
RIiBid6tU0BeKlW/2E3RSK7y0GhTiuJUm2+GVrwQ9mFrLELgcdqeES3BhBEzz4Lh23Qv0vHufPKy
+Ry/FhOTySCw/R4MrSw69o1QK2MP2UeCwKXHLEmnvUj/y6fRVvHH990C6iDB6/IWN1ozAiM2aJAg
GhiU5zUTADBWIidFopQg8/Unwshf5GlRM7lwjGAAeyW/rUKetiNC7kPfW6KqFIaqvj1mk+Xb6q4k
0Jx9pEJBHOZ/Y43r2LYZSdRjlrfUkSNCQxchBwD33YgDzWfi9H/fKUH8iwOVqbfDXy9Qn++Gjkfb
DF0J/Oh9BdUNMOc4R8nXiol0XTjZcAsoJLpVirZZ/Av8PpRChEKPoErAJxzWtDxr2igwc+yZLCTs
fKbApXiGnb2N3khVWlizWwL4YVgL6ky76kRTJoiqIjZJszTEeOeCnRe4LnEoPJ3/ZaBe32hCyUzb
Sfd90QDueEdkDjDatKhuc65q0PFLKr+iIpe+p/GOYGAggnZqHi5meZ9DOW8cdm7TwGnCNflaVqaD
deQK7Xo/Yjzb3YfnscfUMSPwYNhmG5Wb8LMDWfOE4EKEVH/pA87z8Mrzqsxd+xWz2Bj3K+5zwcnn
uFXEEPikWe5KwFS0QG2p/VckAwpQa1zF+humm75oiKJUN/NXnIUjfVBPwiNqPETvxVP7iWga08GE
8ckUVZ9azawrza7t//TKjTbig4prm3DjkvceP0B3sijQp2MyqJYQ24aqrWacF7ZcfdKNoD7cSdrJ
ISzCYUPV0K7B2EIaNjA6U1hWDqEItFPc3rjggvPw/kuYHcMEdmJxsoia02wXCJsQ3cnhNr6Tw26e
xAaaPbLt08PLFdYXzDNobDmI5VVjOWbCePLXgIGiQ7eKERsW3iQbJd3j9LU27nrQPIF0ogRXq6W8
6Jr0fi3VMzgTRzLNKbbh7GdkRxx1qvr4r2lJvQ+8SHXhboUo5BDWa1264T5UOzVRhQlPiQagSL2Z
QFUwsfdpmZZoJxutz9bAy1F1bMbczlwvL0vJ1XnL02k7CzVEsHG3PfmEt3rwKrdDzhpEk1zzo3zZ
lrF1I8RqC/6FqIMWcFBTIUkUqZf+WAyE29g10Jza+MGqrG8Rs24YWDvY+X25wC7hgd4YLv63BibH
Z9JvHhd3A5WRQxpwiER5bJmC5JtT2U8MpP5nRo6FY7yc/bTHNmAobBcta3fBJ9nh6ynmCMKmupxT
FO4619YZEKY9AqQ3rp4kmv10P/A5XMEg3XXBTv8TM3+cczkAedf1AMuzLsSVXk/hM8dyxmoA0PE2
MJRvhGJRG1IqedGDgz0fQlv1rDlAsTYXeSwBIHJyY1awdt2kvbDR6Hf32jjr47MLdGIx9t4k6AOm
HWCzDJt/Czs4gIef4V39gdAYLJF775ZPV65jQ5o3/Ztb+WZpQQSyEJ5OdbQaPx1rQS/2Jk6oitFn
beOTthpO2Gf6kZne1CTDvhoubr092WVe3mX2FKLQVw7hRbEOQaHT6heIlilgCUManOzDTbtW6ObG
IQLhclAkHqIcIDLWkDsudjDkzxHLevBBzXCAwlRJCIVzCd5xtkZ6TE9uXJoP28I7xZr5jSznYfez
i3Xm7jT3GDEBDTuXzEDr/Cc8DqA5UxI7tNSgVh72U3ic+x4sXIHUMGPQSP0gyohS6HJHYu7U3r70
01yZo2vkBjWz8YVqnqjnDhEvXdVDwirtHrWuz9GfxIGpYYUEEOh7zpHqaIsuKtTH0YwsF7L5jHiz
2YRb5/NTQzTB130Ndf2J4P/WzFjhrFHajY6K2bxy/IKn/kszIVCQrRJom2HC0se62Nqdxsd7nrrd
6rNZ70xlgFFEyvje+iPh1YyRkT69B+mXoYIBrlogPEPu1EVIKLQlEsfGsa8Pb+KI/bQrE1ioOO51
tXyVM4f5XjPKISyuUKpr7vHrRM9t6rK4UNMwKac3QGZBCjWyaa6ohPZqkAFWiRkgbZNN5p3AWmMh
Tq38k5qWT42igyQEk9doeMqJsUgwrMbh9V5I8OsmMd40PcPS65vsGpBsFo8A84fGNrQBq2viTR1F
UgvtgH0a8+L77vZsVJoYaYcEZ6M9axcMt6f0y41N2BMj/cEL+bW6Az2Tn2wrZRvdRmxGglMvPurB
jUHuHQtvBJ4ngHKWaEorJInvFoJ9d9G2YEYVoN1I2rGu6btEJhYipmHPYAG8AYzLjD8VecJwchjo
aO9OYzFqcI3ckj7dsYotQF9+SBY7bhdH2knkWPkbTMVfg5OM9RnCKFWhTZLZ8gQdPYQRIxvesRar
VoX2hukg0fYvRxe2oNp8ij6de7mU139FOIatF84x4CNz87Ra+ezzxxqDYrFmfIULrZk6gh+V2xAr
VOCNmZ8L92NlOFQpvSefC7qgOBi0O+8PkSTwKd98mNOvJG9yDpkO/ZuGoKcvUbbqGPFTqFJm7P07
shIkFluodWH5BKznPapeu0eBgElsu2pKxI5SNJTDzILLKyvQ5N5EkuuvNYZCTioSFOWTNqWXOEtw
DnxIfBLjZsgnksQa13swJfHBqzkF5ZaZi+Bf5yK4l+W7fRBrgkNGtSNrJFLOFN9AKWqg376ZyFAt
XiAg62oxeOO/gfwvIdzRILbOSmJVhxS2HOJX/O7/rNiTcyxvhghSbpyie/BEmpsvBJu5TroF6riH
YxPdUByetPAJohySoLHnLo7OyXL2UNQp6hF1RKRAzU60SNuLEchb9fpD3sLm7DToTEP/548SMcho
3I5PX2vGfngZyEKftIERsISqsLzaMy+KKluC9/eR/Kx9oLowV4Bh+xl6+EPUOaSxVZ42Ql14hwmY
TjAJ+pf3dE3vY0KV6/wDrxXECnhB4WgodIldAINi+TGtU+wQClzjeDRr4eRgtQtf/BHiYdkfC1AK
Ru3Qba5TlRRED3LYBDNPwwaZS9LNIhnGdjmt+zZVEW0T8wpZgk20CA2MmYzpz3LspLRSHuNF9UOd
QhebiHeYiv0jW900mzZ0UeCFBhDIfXJzwAb3MKEadmpOqrHRB4/ECg/S6ws60AjAOfslcAPqpwJz
+cNlyMVuxzghO9lEtcCZSbSJzT/zf3M24vG+qD0jtPk8GtFDh4qT2ou+XyqAMi8ZnQWEpVbESv39
nRZaNci7OkMK+Uxbg/mI4wmmWnZGtzjks93HuLSO0jDcjxFz8AuBiLIjCZ1m7DBM3+X8U97j0J5S
BxS0i3c+aGsgX41VpYwuKqsnNYkgP9GCFD9T1Zq5nvyPwdux7GI4nd0X9Hk/xSZmmr0hOTsmg/iv
KNGTPu/51zLCRqCdu/8Fc2lGxmZrH01mKtXHhdZZrwukCnvL83w4B+F/Kdqz0/l53cj9o/Z4s2hF
nisOciqyruOMV3jJcfFvU4HPBcS96BGbyoefus+cBwlgDpL1hGbD1q0t57C7+9w2dU5CFOKCFydP
AiRSYhmikeBTc5tAuxx9VUyKgZ0/aUiP/IyQQJd/us5nD/n5bPD9R+YmV91M0YF659JZDIBR2eIB
hloH9+VulWJ6ZQYD0WDJ6YvlsXeTvvSQlvu/ApmzUTJpLevwdpS5F41IQszo+PKe2+zBgMlUbgPb
3SHHJhA+UTFLqCHyb1gqNvk2ukdtfuN7pGEsOrjhcZRXmS5tn/eJ+0tfiHPhZVMGp4ixNXKQb2mn
Gzx9WXPE98Eb2n+TpfxVMdOXATGwys6Z/56G8vkK+M8XXGlFzxGFC3k0aP05GWr6l5svDNYgXgnk
N7i/Pl2pyGnd0rkj+k8OjQusLiNYup+IlRMnlR18tU4KkAvtPnfs4s67Qu1kgb2jBHbKsh0MvFj+
sebM3sXymJ8fG29JDlmxZTfOY4zu84MvzlNy50TyzpfHOh7Jm0yXONoXSmObetb1ZR3woIwf1gfB
bFr40EpGpdGtufjn1VY9/Cg4yVIMni6f3d6+yuvsQpfaGgff7c8pk1MRdX8DBS48pKFUGyk+cIGI
4Oov2F5AACZrPOwOR+Z2nQMHWp5j3NelfCT606hNjSE/fvKmCeZuKhvpCZDHsjWmInkkIBdenLk0
drn/GPaq+DjLnA0uZhiiD3HTlT1qDn98JQcpgfBF2Gff+5jzPb+QonMZu/dK2kYe/m97DSHQcxnL
Aurgw03NTyzWl2vOecOJ54eCk/G++2vFju3rJRQyrOhoVs564d6d/EOud+966UodcPoEDHCTC1qv
/njJEWXb2e0cije1Auq2GmClRmt4ASe9Mefxk76QrnRp4EaZoO+WaOyw7KkgSD2x2kG/Nd7qAZB2
1uueWSogt9Y8mt3nK9CTSgwpze+LSNOywcqtXMIeIC/jDMMbVW/jzsATqrHDQOJyDjG5v/9WKfL3
2iE9TYFhJXQk8kH59QM2QcjFmuV/113/Q2X2Zq6NEdLXoPQVfreDG0VfVH96IpU+4Hni4uvNsXm5
1BObdDtHBtRDF04zyHqc4URXDhGlA7cpwuWYEOzDV2ltqqKy+RW5Nfgjm3aZ3iKaY8C4vF8dYobx
TmCK/Jw9yKh/vkFzKtc4H3nzmvR/Dw1UumwbskWtrO6e/zfmEAKAEJKzpJiReO8LbFfjEODJAVIL
bJ19dnYL5w6w6MeV07iCWbc4x+5yvRB7keS/Ivw2qgJ85DgbacekanSJ0Zl01eMlDkUcXkR0dLXF
n5y73tElg67ELZULKUDa+mvE7pqJnv/3VvOjXIxeRjII4J8yMcQQEiFx7Qr8xvi1eN77iokBDf/8
1fYoZWEGWNP0wYJUwoQOimG+RYyTotpTjQPAdorPE/B2YecwLkOpdIKyqAxf5vnRiIJ01Fk+REkj
Zq8w3GKXFAZO56pBUIsJIbzxK2bcaWqygeu4qYbVCdClAkKTpXcr/u5g+KZdDrofw+BdPEzbxa9m
7VFPbtORxRl0ajtIECR1H1NtlncSMzuwmU3PjbB9e0mGIceoZM5mt2T4Ez+XW1Z6UQu39qRSXHCz
4Iy5WyvGBHzimQQTvuq+UnyEutdgvi+b6Ir6AzhRyrmfmnzObJ1EF+cgOZ91WYFQB14f41Aszboz
/UnW+xFgKPH7g830jr8yQewb4M66RS2ptWRlLCgYf5q1HfxYTO0DKC7b9GvKOU+WTLG55rbhmMgJ
8Whc7CgRfma2aNQ11QuN1QO91I4aS2oLdIAtSeW5J6ye+R9Qlb4eKsg4YVMHVpor/RcUUjprRk7x
gBxQk6mQXajExjpY4yKJfAvdfp0c/EZfi7WCsXOGHotbi7/XjpSg2OoMweQOJiSGbcpHiAZSOpl7
3hhaeWB4FP8DyBuBNbv7nWiKpNTj69OEBLlZGVZPdphNqdJC0TPjhNl4WlWOJLp/VDBEeh6QgoNX
WmkVUDJtfyEC/dl5fGzzoHqgTz4dwhG5HR91k1idTJDf+4J5tDAwzXFC7wotwfNgRDB3KP7pofdT
DN50Sm7xzNV0uCBPUDGjAbKOpTmhaWGVtGsbC6pA9ZdjQIQRrkYeiNET3OyXz/xl3+W7gwC8qnaV
7ExvPShHPQxwBoWKKiNb39qmPiHWFKY5Or36sfnwQQFztwgtldKjgPU/dcHFQGLOeooflOXlWGxk
3XqwC3G5tNO1yuaTAMFrZdM2lO4WM7f8q20O6tHAkr9D52+Iq1kb2w7Qv5cgo26kScwfpjIJL/qD
yIMG2cddeXVu2DfQbamPsvYzego6Pk9L8aOGOMe4U0Axm8N4120klogI2ocMleZ1Ql+XFqTiY8fV
7Qdf4VR2R+3prXpNPg4LSIvJEsZnt5orD7Z1OgzlBHyzaSMmV3SPSx/BrbKDm0H5z8Sff1Y3mBdA
kgMCIjlbGTuRpTkqCt3ADLCvT8QnpiAEgEprWJtcphj7vP6VGV41JJQLK0R2HMlz5X/aZLg+O0fX
T5/cRn5u99o1Tec1mB8zDcljzLHyTivDTMBEAz+QPA+93irYOPcOSJZnYwbboOl4XYJDG4hhxek7
DWLfhmAH/MuwU+PlCf9VEbXkeqnuFIR0GUxM/GisTj4wOPgZd491ZmpyWvPyoGxtyLrjwRRiHwmk
G1zqsQbO8HYxq3/Qnvv9afSTOGOm1gk09JggKhIBtSf+7B/SANUilBDwrhKJbBxCHWJSvRYbPsns
uFhkhpszAybxDow2vjfS/Qtbmwj/jmB89xf0lRvpNL62pwXamZIwxVd4v4ZcV5Dkv+ZtIzr2E5ik
T7UQI3osLUgiD7AXRWc904c6SAngVMAFkWkwt4PU2CyQDjgT6GJOHbCnMZg4l96Zi4638kO/Cqko
bI0FBrHc0HvODGfJTLsuN2d2VdOPPnW93962jDsDA3UZ1Sy2ceVHO8F0lce4m3p5PDsUp84AhsJR
QhOehzEeq/qP7AD1UimnyflaMmPCw5AcW0N3fIruQqUZ0LC2qEImisDhfdK23qOrks6aQ/jVr+W5
QuMUSL537UnRre3McZ0YkfcsdHseAwmGyTYp4kCd1Npx657ivV2alBQ5P4ZdrV1eoUNx7Ufo0EQl
fx6ILglJEvassb1ws8XLIjNmsBvbG/448BBq80uxqxbXYWIImH3F8P4qRxBRUQZnBiPD2q+EF6EN
uBQ7w1B2MRp9kY1QETPykA7ft6KcVaD6g/q+/P6iBzFPOZlbmN9qclOH4aGWdDXXwQkZpjpkOBf1
RuqM/ElbbAG9yGf1ZnXpy52mPebEndqOTxuWFgSFAj1OZi8PA2CZB7DgDq1vyAQlszOP9iNKw7c/
M3JUalfKV6mb7pox5/CGxBEFXZxe7C9wJkixhTjRi0mhheAnyVyFItXVMgKIee+ndZ08gfeB4lZa
pWsy+Kka+36AavZitCMFMVRT1h6t4Xl0XMb4cjTWe1t9MksJyo3lXd/MptDoIH5fCmN3jYm3YYgp
gTQ1QpVfkjFf/0Weu0eWtYY1LpQl6RAxs1gN5n878WSgbrmPnubfV/ynYn1MPK46Zv/5LsVHkGme
Js0Ouh12o/1BFuoNSOpus6sK7S4+JUK8cnXr93IO8aPk6pLycT0lY058rFvQ8A5L6w0Wl0rsTFvz
0lxJ+CBsBrhecySxYCR+RShPIEyE3gfmepWiivezuxI6/K+h8e6+fk3TxFymfuVU228f/typLFft
oWDTI/enP9v3oHIXhSB7nvL6FU7Gb/8zKp+bsSE+fDFjofo5yuVn3eD6E5fsicSL/PtQNYjLi5bQ
egn8Zuwe0pGqtU740YKz51eKoZI8PWMZ86R+AUxEWeksKoo9lWZuyX17FJsfcU2L+BWGaXBseM1j
aCjRvvXKkcQFdwm3nkLBPl0O3GyxSmmrZ5yCwtO3yOaCGY3ygv+Djev738HlYRUwch11Z6ma6/NV
OfyoxzokrOLjV9cKN2kWkiUq1ATi56YgFFlAdT6iMWb2v8PZnZgewZoH/p06qn/9l4F/qQHVz9WO
BcII/MUNSGBOW+hEGdmHE6CW0TPXQYdgXBgyEzI8yFL2MFNVI19wavwuq/O9ROvYa7FgpKvAmVBK
TT2C5aEkmA7VVp5vc5+7772icuauPKcRM1GoDH/8ZlzD/65UFhqEhc4mXS1FtwcM8aL1bHFHwDcO
xASREflEcqz88X0Wt5JUQxitAVEQ0Ceu/662TKcr1bgbxy9wHKvVDXtU1Yt+1CbbFKpoXDTd0mTj
B22G1uSVSRHAwuzwcHwkh6xJNB/q3R+E48H/JHsHJ8wpLM9Bo0D5BI/8gPYB2ELcQUIynykaPF+K
b7J8OD8phWc7spGTydHqaXirARCYPZVyjT0iPTFSXKbUnSqBtop5JK3MgCxMxqKeMq77iioDMRGx
+2dgqD9Hxb66TPFYT50kU9xfuysarRW48DBJkL32nPm6bPj8LLv3JRHhrw/0G6Vmlkc3hJEZ4jW6
PY0f3qoeVsQNh3U6coJ203rErkUahB8dSVgWHpNDPf0l5uQ0QWSkJV4RSufXdkm2kc4WcJXU9uUK
Gi8t9FuuSZ+xtlKs/8ycDvwuFFiSlBLKnNPJLJ3A7JIrRd8ZmRU2E5E/n7jemDmDAuK38c+RvSxL
zou29zTnQYxkcSPzdJLK/jLZIOOIIBfj5iFxCnJn5RXcjpTeas1Sv/5T8YVREs7Ajhh0tgaAVSMt
3646aIcLaVlnQcBY0XO4bR6aq+TuVorsBcDS0A1n2amRXjRo/dwIqQkGAQn56bM+FBFX+25zLvOj
bVSHy67ZKAARTbdNye/3AmVFELGp8nLvQT+3PFxKHUNu+BRBPpsjNhmQDrOIf252zSX7CcBhpJsG
bbYR3TFQcOE7jlZwTzOr1kd28Uh1Au3Htd4SSc0nNQh6F14/WYmt4yk0ZSJ52F7Spg+8VWl1Ow6z
AALH5ZS6RF3CJgTEoR8TSm5qDKztsfleI18g8zA0oJ/ZKwSxfkqPZrEdwdKn4+JLsqfcDWAlUmKV
zYigM04je6ZANOO+TgC6+tQ1HqZPxAsvTVPYoDCjihNAEwGJuRk7CXD6+75Bnn8pZ5ueZHlOfDCF
oJzs15SPezkpSzaSxvc0s1vVnKcHtSSOZPtrCqSs7iHZLUCib3pIDft0mfpd+13qTV/2RcfNIZs0
j+YQU0OErs9GY6vlV7/v15YfRO/KJ9n5L5HnENrs2JMBh4nGZdFMj1thOtjeZu3R3D6GQ4TBEftY
9Gw5chSpJeuwuidfdfI0be8fw8ObJ/wbX7PZ8QZ+FVluGFq2+a5bDeA2scLmS2LG/PdE3Oy1AR46
eIwfp9eTEwZaIg2lNwWOHvylkjKVP0ElfTr2bOUnJIQiAydSi+O5DMLG620/f+1jBTrM5XpM3gmD
RGIsbBsgyaDYC0OV/sQHGXsnQ/u9ky42gFr8hh65PtzPfverAE8d5Xxry0i09WUOAkMOso0jwwDJ
NeENDvv+7qxqCvD9XmpLsxQAR+3SeKNmXpi+YMRVjMDtNnos3WNY5v51YGSPKAYyvg8Vsgg3DfFJ
49YbX38ZVzixXqVdfKAMU8dxqyZgbPVmvmbn+9dJiUp7nHF12XVwFsd5PO+oU9IMiZbusqzpkypa
Tg3YRdoFCP3UoaSTkTvHqg6rc6aUB0Qk9sXr+xo4/GUQDe9vqOGHEv4GhtQncoJhA5G7nunNDIRU
tKxbvFE4ecmcP4YBSebG3+rMHaaouO/+JmbR5GsnDsfP2JtTgwCGAK7vw/+bW0MBVz8G/h7nI6hW
Wf8xHtbGVU//NNcmWl/OUIECMlfVq/dPjIKFEh388AureFllUTOT66zbuAipWLIUVtE8YDWIe2TW
nFJXx1RKBgk4f49CIc6tqKV4QWO/LpdbawWG7CtItxKXLps1NcAa0TfsVFL8PS8cXnkw1pWs4+pM
cHK+sH/J2lBCQrtPOT5/Dr9ph2FugFz8c/XW1fCjdBE8BmvjOvjL/qIwrwH97tdvEhPqu2SJ0Qon
pkt6k/OBcNstS1Q4n/q4i1Ffe946zpty7ZvnnjjWt761ij1oLnqCloB1cBqw1UdVkB1uLn1Cj2g/
7ucXaPC9Ky0elgwN/v0dS8YgE25xIKL32LuWtPon40E/lk5shyNH0jZY5SzBZabhpdJxSFwmqvVO
wsMlxycHNSL6ghn8YCj8ghdWQrBJc13VOqFwUx44tUSBWwWtj5HhhFXHfKGDxQwMv2s25w2z9elI
fySVV3ZE/Ln5afUyccn2C5x1OOLNkilLVih8mzthPGxjuHz9stvZ/747/LdJ1ksv2XHSry0UPxwR
oWEFyl7wJdMJCvfjSyXQ12AioQskdHBr5wACrGdhmF2MIzj/06xIYsCxZ1x2fmkbOs+v3t7gFvaK
93FVGjtPJTvV2e3EyBcQDbSOi45qh1hfHId9k2l0exMhWLf5dsqQA5tKaAQM5o1dEN9ao4R84vYf
UjKz66kMa66ugfOokTP0J7NR4qxc7Y5z/0tEcSbO09VAGdfj4INPiJpxzpaIFXred133OT4s4+7L
CGAvN/YQO713fEYex1uHj+mwlPGibKKWFcV2nz7iLMHQS7R7NP7W00r3KP3GgBRrdiVmb5nW+Wau
D2LVMJyxXlpY4G/CExqCD0bJeupPNKq7O2nJlISvqfTfcdXyWTI3UilBaV1foaSdPVIuqEAuO4Si
MtKufTelE/WPCh+roVJrBrHpcz06ffpAbJHjYiLdex+22nkhnCd76ueHyoR2r3Ltl23BN1gikw2L
7F1SIiIBAnnijgeymoIXh6s6kbTlS9pcZ1udQke87lTPEeVX0czKgEzddM0Q1SEinlmeIV9PpSlO
5ZFX5a1ssL6VR5boJNMm53/8s2ScRXnbodYk4HIeAn1uBKl7HVQmkQllG2GJz2rUaBom3VTeUnRQ
HS3SkKlMNzTgRjjZjDfyM+4Y7kgVfr2xviy35m+QItjq9SJYJHQrou5NmdfFGjbA2n0EQnFlmzFb
r/Ll3oGgm+vlbxjZWLA8ZKqDBgWaP75/8EI/nDMdGSv77tUCCbwbU8spnGejg05/jR4MMYTvYnWx
W61/DAgVvUgYYGLDbyzC89Sc+qZ32VJ4hWLVMI6SfK2aSgrFsJGvqXMk1GCv2TeeYYm5KJLhAhIP
41XIiKAJEraErMngl40vJdE+cmP9Jo2qK3o4xyfI8S8tNrnBxdIm9KgvgYPkBymIrlte8hFJJTZr
rxEd2zVyayO3H8sMpMqvgbDIBdHB06MsyWiT7AWrzvXBGQwyr24mqrmxFJ1MxCzWydQMhAsRCAAq
d04IuQSFCRdZFz5ykpFnuDBGW86+UfXr8bfwz1BNZNNsTBIuvda2opGhs9lzMhxIbZV6+bTPqrLW
p8tVyUKts6F+Pl25NlCFCdLTQxAzwNpDIdFCuHG8uPuEMJsfTCicC3r+uTMdZ8Pm3/oRxxOrH1mp
3d+bnLY6fl3MQqdNH4uG+ELY5yCzBzrXWq/K1SL+OOLoHCeom90X0UStTaPaSGh+TM6719Stj3Xp
F4Vb2z8j+yDJHT6okrHZsA3B+kqqbZgg3D6LTjY7qE20pbXr/hs+SkPwCBq7xDGgcDURuSSRU61h
I6skbgz4ZSWESc0swIWyH8RJFTeIE8VK18gt/hJzGIYffTDJAe3dFOmVPPgmLtTodxWgKH0oxK5p
g4WBntuHIyMz8WpeQd7sAKxpMQQddrT5NUQcIbBav/m266lldoXsCpyYjaFSvh4InbW7AbzBkOQ3
edz11yYxHgF8FovKyizJm+0kTaZt0foCEuSshE0og6xZN64BUc0SdZyeg+ghiLd2O7oMPBOFb6fF
VfnnMvg4zj1Fg0vO3s16KZjPqXBQFzqqv10CMiSa9/ZrksdUUad6LwShnD9ecVhKnl02niVqykzV
HF3PRXvq3/CPNHPcoIW6/QvWwu7eJxmGpB0GgguYWMN0gwCIgdznrCVN9Lb4Hd1HGhSKzKcMA8se
zanCCX/wZClLw6t6MwmcKa+V2xRle+mdWGRVJZMu6mQVqZazTBkjB/1Vz3x6IINmJhdI+g7hM6HK
DYsAirKuSuV8XjKU8P9dav0idiLzr7ImGHxA3ZCD1zzHihdhtyeajJFSmjZg2Vw/q3O6Fc3hNBb2
kcLXpT55TuTjbKVt6Yd8t1uBzd8ntJAzii9wEV6GdTn+MAqhlU6k8D7bq2BzBfoe/5l4hXYikw7n
Tj9nxNw9O4rchFxdxc2CAYk9/XMVtOS845fD4DKxE9KiBc8QQrQjH7jEcEaY5cShSLKjiP8+Wjef
kNFKyK/386alPY7WzgWr+N1Iu0l+pj3rO4qTP/bMkzKjgSlBKu2Qv4hrFSUGSiAWB9++iZ8T//7B
hYnAyJjuLqh37Qll0cPBT4NKwpOJVb+3hIWjxzAdkSgG1nFYFaO8ASdjQmmsY9lTkG5VKO89K4B4
ljEKLh9Ibc4EdSv7wQVvigra3YmnDoKY4sWIUlJ+d1gAXxLYbL1ue0zrQg8n47cMMMkLOm/We+4o
yImXUNpLxK1U5elok+gRWTua0x3kD4YdShD/R5C3uaLdEHHJzP/b7fMRl4RfdTDR+4WuTs2n/E2v
iGPuprQt6sf0D4/ZAxEeKwp0OY1OcoXvoYkF7vjGZ/jUEraP8Samlj+D/H8Bz6HRFdawvCxlmInd
+eKNkSninlaDQjZpV5vi3eGK97paRAkF9/5S+O3mLR+/icXBUVBFbzuQpdSvAVVFLaB0kmTFF6qH
PWkusqU/39sesYHO6MYAYISZ1kBRbmsgPYa4EIJu8+tJuzPJNOacKH9tp09attrW31fTMvfJMfAv
sDBFAnzYBb8ufReOECVS0rlaW3Ys7zfTTJcwWUzbkNSwaygUz82TWNm67g95rBuwZsCRhoNU9mU8
RN85Mph3QMP7OA/vYt/Fh2zeD09stRP5tWHmFuvCPlrM+6bQMY4b2Fjlu+76Hs5xJ4fFqbOmfhc4
Z2mKxcVXxmopKHiNZuEcl4l5grKNWpjDrv96+t8l2HyAFWlwXLSukrQK7aXDuvCp8rPsYZ5rvAtR
srg7GUCjpe9fSBPRPGPHPz79G+86YK9h0KU8XM65VMWiBSx6wR1q2K3xD/vFo7YPGT05VKFVby+b
tBIl9B43rVt30gRbjjqI9AQ7y/2L9PKK2wF7qP6B10FjeyhboRWrXz4Q3ShnibBpZVpk2LavjbxR
63WfFEfV0yYCp+ULkNdM3BbUgaEi2AZphfUi4rg6TrSn15aWPzk6wpfSxp0pmSVu9v8s0Bt5Ud1U
Dd5yko0IAcQOxImTnrZj4FDUFaS1euFQDYLnuOX2FtjR0GrN2EOztkeZg1lZUQZfcPQO6Kx97+0K
49F9S1vJuWMytim/lV6oX/HGwpfFMenRT16C/aT206XQAKMTt8QcdDlL8RLKa0BsIzWFNJmcv2W+
Z7fe3nYBDDV9asE1uIlProm5BVhDCPK77QUSsJhXPHiRz5DNYT6x1Mavl+PayLnL4CwEZxGfg+u1
R6Zzc/r+H3fYHXq2Aw5e7Ii+dePAD1Ae9LJW9ktJvB7lPPIs+hUIELb9FZEb5+W4bE+jDHNAUMo2
gsWNal+HcXoe9wrroPSfLxeMFbIr9yvoSqHZnQ0TogrG89yXh346Tsg6QHWxt+znkyyAjk6jyCeo
97M2oImG0m3OZvWC3Dsu04PVhS2GImch7YmigaTusC4GEnCoZILoGYRoRlAb0uacCgk4+/xNTkKk
lt7Dk4pUq2tTv0D8eXMTGT56NVR3/t+dzVMhUG4PzFPplsVt/eAWVxCZ8i/JBW8z4pXh66Jk74Wi
HE92MTcztgL4W/LxB6gq/7CrvD7/vcKuXbR4HQrwAgH97xIk9ZMB3ggwRPhoAkal9H/537GNkvhi
bX8vL7rQZevcpCI18WxQABwSSJlewxi87VwWr1XFGXaBxVjOrT9d+z/X9xXPPI5fmIOfhB4h69gg
ugS0NjS5AI6X3zB3bGAGzxRMhUXSswCHlKvxsCM5sDS3y36t9uHVH1o01F+KmTos7t5nB4dxFFb9
I1zf/Hr7sjZQld1tpCkjlmqR2+nQ6RULphwEQzsPe1FDWHjD4AWurYaurPMM83hNFOR3nPkm6bdU
2z6r2Yu26Gwhs0MxKsJhbwIV9bERQzsF+QtjxidTqbQdgYKlU+wfYNeCgla3ly5nkSn0AayI2bcl
VFNsGVvAYKqk9OEJZcaGlkC1I1h9zlJUBd1m1nO1e98d1gVFUHctxcQT2wVpSn8KXsANPFl0vO9H
w4l0N9g+x6Vu/kNfgQEz5q/s+iw23qKt9CNgf+jDKWiMYHxJhkw0q9wKad7lQA6iqQ/veur500g9
fTgHpRBw8xY7wbBSJHmH58a3IWBu71K1gCV4BAqB83mzZOXlFTjnIkIjt8SqwkZgasHvj6AaE2bg
/RJfxepOo9Oc7t/9F0eREXUyfDDJPgIHWkuYsy82BbRtA3v1MZ+kId7hfR7/uQO7MtgPV7yDrNCU
P/WrTmikbihwEeby30I1NhIoCF35upDCdv1W8Bn/hlxdFR2VD3+S8xNSdA/9WfYdac348KtKj36b
F7P8CiXHjrv50t7UGG8FDcxc3of+MKSsYlF1TTbSrpcEi2SW9xGHl2Eckel75QH3ryzg6c6Vb7eO
Ee6co/bG3L1vFwdvcQkkQ2ncNIhHaZEbEpNRYrk/YWeUYuatAmLx2424ApOFMBzuP2EqrnVRdm1N
OPZ3aRizxfLtEoXE5MBzAY26ALCab2q4/3TwP21INkvCcYY1oE6+OOzlZZRSQaPfz2SXJafDpAdm
C4spwh2N/KczdcN/FW2bcU0Up8PrQG6+/7YhkLw88QxHTXoT2vSo0UwXLt7glCbIfJ6TkbNwkero
oQ3wRwmtF+/L2wtQ10DR2u8o4pHDC1iNmlXidmgTO6kp9sxSCuE9jOwMC9vy1ONFXMAut44FkxNI
mPfSP49vwQFSXWr4MCld2hDD9gNduEYOrbx+o1ry3R9Jbf5RSWC5/Bz+lT/RVM1b2hZKS5/g2YhU
IaCHM2uZy8tW7KBMeLRJ/F8R+IWIeH2xGAA60lTvv7rUAqlPnsTUOWZEmXgQWkGzHaqwq9q1urHs
tbcJ+UodEC1sSR0QJKP1K84+uz7eY3ty9fBNMIErjmfOVMR9NRChoKsuE0z2G0YFBiMuSZlyXTbp
0Og0kJkpwwTqBpq3+qzOwVXf9fuLJlLxiKYBg6Xh/eO45EOtw8F/d5UGUD6lNhWj+qTow/5YyBNJ
Obz2vGK0RjLikP6US6TR9dbD3rz8Q/YNj66ojA7008ONQ12gMw8ukZhfBKmq7AHIlTF4uwA2wjoR
EEnbwQm8yoA8nOYd/AfQagrsu4fv5c1p2KMkonOUzXWBMKUTD9TRdxmINO6A2iw6ltS7DarkOlg+
w5RWXlXWJmKyT8YoFNLg4irLn0aPdcRzGEx/CW29KBFrGz0pe3mTmOojfdlg+YIXmCkozMsqKrFb
G6Yaq6MoocpF5NJuV2Cdd0cOYnUKlq+VkzNu3/FrBqFXGWlaetzebwVV9qhw8eTnV3ZGTJkygstn
gUkC3h6MK2PelwMrwvKL1V+uEREkQ2LbiN1IuzbyhImOL2ynKrInLTo6qW74+rXEOdHZOy49U3e6
Yka9kOJZ8VVoljf/knnc4CTv9vsES6fZ0jyAu+YWnjwQzsl4j8KMD2H/m7zpn8MBsEUTIXEArxK6
Sx2RylvTzOb3XW0qMGg5fp4FenKxcaHdPsFY7od/YiFlpv0hvqQQ0cI55rg0ZUFcpamxjPgeGJ3u
q4pNpBrw3kHSiSWqCw5OnJQ89FrUHCGeY94CcSmrDbSx0IUsX46iMqwsPQygN/y0gxYeQtlXd8Y0
YQ6QK9CSysNFY+QbwP1TgsTw5lo8JORzZAoHDOqiP/FuZIbwqAcx4f3rzKbaIv7yNi5NHTdhyUiY
kqMfy/AqGps8SJCpFBizwbnjlt9+oPRlH0GpkawNiOw0mAVIsHxpWoR8IugNpELfyjoJjUmaRVhP
kthvGDeOW421/DHB2Xr2msCpeuGcFAKO8H2l3bqfK6OlgsjnY/yR9b3DC086te4IKHFSZ1+y1i7e
tXoPqQFnevy8VfuVQXE9IPIwMkDmv2ncL7QG5I79H8evZV1PBbOjaegLr3dkwRQN+VtFfBiKVRSN
goP1IAipITTHsgdz15QgKZH9QaoXL6vlF0phyiZXmL6RTNLUDBfiNpSfbgo2Uaf1a59HV8eTcDBF
PLzDujkTHBHA2SLVYOHrNSpwbF5eqOrbJHG27s3UZBG+80Hfa3X69RPPpjVgEgZi52hpZ0h7Bpc3
pVWRUBOhhzVo4W8/BlRCu1ggxtF+FJVMa7NcY2UvWu4Z89QlkAsaxINTShSK4T8FJP65vbuPyyfK
fWOcyw2yhPEwzg+gLZTMA1novGJIBj+Umzi/RVo5r/FBhCYBtMv/wW9jhN6dUYUjIOdyq4O0mGyn
+OZN1+AmSFZlOAyLc/9ZO4U9vEj9dzkybnAckGwU9teO1FWrTV4XyOFh9613PdvB0QvUylaSrLrP
uD72fU0VRJa8WE0obzs5TiwAN4TD7Vay+w/HQeoCd60p6oARMusaIa1/120OBFZBqmWYV1lbm2N7
EjXdkXcFZOpKQVBkT3pxnRTGrgIbZE2OlUu3cUln5+DL3KgVI5bQZSuOJlUNc4BhBXOvABYJYcQV
80dCLA1RzT7giRjkISNkuqnWTTfBQQ3DhSiRVxsx3rF1A654nluR87RbFQPvA+qci/pqQAR+KMSR
S4dvkrAUUMmVolFM0bv5hgsCKfwmPZsE79RjW/oTDbUO4f0S+nQ8C3GUrSkBEsSr14zVcy/5ptVn
DkNi1iEntu8apIUVakpvXegP2KwWwtIxw8eRZJFw0EFuQCddJux6TXB2tY/jjZL7BBeuYGj60Y4S
Dv5nznPXxoya6l8iyvxDTwnlsIV5sUsjkFYvDYDjbldDSl4B2CtmBe+Av8Ff16nKQ+0cXdlDPPH3
QojYITb+xGoWAxqQt86EHLvbGsBjIN5UVI27GrW1Zd1M7C39L9nZqYmDXfP3YqqVR3amKMMPVddN
9ZHheXGN8Q1aoM5H1PfF3CIaCFmvP6Rdge4S/vovUzecPNA3OuUCQVmTvBVL+tZROxYh5whpPZ3E
+0vvC4Iky2EQBoJJxgS1poXY/lxpk7SDfZGJ7lIVIMvlDzpoS50KD3kNiOn8eQBi+6h047cztq4L
X7+/3RLkIJqpkibUdsK8s8tKsTZyogB4a1NN4Gc2sF86lpLxxNI0BzS063/Zww2nMKV0VgSP7m9W
4IVz2hHCyeTB2BCEmBzxfrGG7dWMCB5B3/69bRApgLK7By9/qPm+jq9mNA7gG4MscSu6frn3IXuR
zf7bwgBU0JbwORDqqwADjse1q8baVJxAgmdJWf9vTg8PLCmUw2iQECA7jayvOxxU/1lggUXBTbnF
5LueN6+p84YPpeNZ1t95P2QfL3zOYJkgws0nTu6EtxCdOFX2+lyLMqc6i6TkiD42dPrf147FkfBw
n6SU3DYyFD3MjAk+xGY/T2plk8kLx9NMmTLhUB+B16LJKVXGpf20jmBhfXkKfbDw3QkblbLR/F/a
gTRztUsXJSYg0gXVmWBZ2YBMGS21ShfVNj7Ilyhi/1XQGT0CQrRgqqy2NJJ4qaKmloqcpnVgKRe2
wd6g1/yE6S19cOHo3ddUjbjqiW3P326ybkEifIWS2uGYoPeSfIX562NGIly206mFm7n1DbGcKF2X
NSCvjpGlgijNZAVanbVJnV1vAuUZmawDskF/TyoTh8e7PCdkd6+jPcqDQLu0bgkswCF2VklmkGLt
P+eOeCIRZSZ5HdAyNhhlMPO/5ERof3zJbnXKXgQqronsyo22W5CYogeL0M/vEPhA4b3l75tYKNRz
LDoH68rtAGQZiY73WA3V2rHdFRWRURCcYilM6JvLlhEd5uCbIM2Rwjj2UNxwAS/fA5mfZVORL362
Hf77jWquUrxWeP0HDLOl3oGHhRnT5mupQJu7nnzbt3Q8j/JTIpOCAyVbelcNEdSP1Y8u3bKsxRWa
Ntc452mkV2dZ8RtNmUmFNrZtn7HboKdDyAZQbPZSrv1iTkYNQIyZSB2dxjOEjyr/utFi4SGieie5
lsfuR4UtS5Ef+Z0ZXxoUSdGIpmpxqh1Ef2orA8Mt6oQz21+KuPrVAgLIY0yoAWt1bPqAP5Fmp2bX
3eB+xHkg6ZVBG0OwS+CWKV1E+JRCxnMUKILmWVfNIBDHHjQXxElgIX+Phn6QuGpppY3niuqZA3Sr
zPcwFi9YSVx4IXxsQt+NY+zHXIM/z/3bLOS+3IYTgFV4muiwjJGWgjgokMJAi6a3IIDfY/Mx4f++
A30gWz6+U5q17hF0QBEoaJU8vLuyVNhuRfCiESlSjOFMbpnJT8e1MnMf1p5qnqkK3HWrMHtfq3D/
umic5kr+EzXy/tvv/cDcuzU6FrgFnzrYz0A8+LH0wt5hAd++oSxwvWIjgyQduI2YGqYeCMVft21I
e4qukAUR1nFHjqw2qK5+m+JdPPWsnNVDJHw0msfl9ld1CdNbvUhpnmGB/51a2G5vsoJ3ssXIc38G
PUPc1dPT7MbxrvqWyPdVQ0DJXoJ8l1pkEJQXHMQPrMVxDejkhzDi+htt0qjdEIqwN7whMizHZSmo
uoKWtMIvbT/goePVeoaVqmtjtJppC04aH5rJUg+f2DCYnuaINSU2FPgWSDutgI/nl2fve4gEWdbE
fX1hznx4kvjcKhkyFVtxYMLGGaHyZIkCGrijph+KYPb1jnJINgsLugjHZ0sxK8iGtiBU5fCNn1xz
m/tXXOmd/NioPly2+qo65VBREwv1av9AgQ2Oziy/wEhY9oT35cKPFQDBBt13OIBrUUupXrBIhVkV
lqH0UsOANcIeqfoHrg3yyt4ZUgTPqzwYzbUzEfz0iuaeiMd2waT2GpW9X7Mv7Z5Tvd5On9YPIygH
21uykq2JLFNuHRjEEHrcJPn2ra2CWTwtVdU5x2wMMtSPmVfynEtuNeHEn/3yHmPjCO2w+kQWk5Ot
oCCydvM25fW0twlIoiycfds7ueFamElYRG2qLFEPvz+xfrQ/zPogJJa6cfUXomxwSh7Oha4klCyH
w7rsDAOh34n7ZQlSkYlF05WjPdp6MaLhUcQ/NWLXcuraDMeod7ayiVPtkGICd5eapA1IYraQMvSS
h7r386uaSP3haeSLZF8kvoHqBnsPsZi1c3G/QgB8pXNcr1B1SfGHESqe0Oz0GHyYYYuxFsIwTi19
GspJONDf1yKoVCt0lsk0cl0V8aiU1vrcwzbGT1AiESLNPfccG0Gxwq6VjaEwnXgbVd2TmaGiZv9s
qoEs9aM1jmzs1W8T4N2ASfZtS5ZZ3ntdUGjT9a0Q0XqJhga1BsByPOMfP/pza94Y9+K2Dsbg0+hD
C8YSy8Zd7o27
`pragma protect end_protected
