// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ypWj67kn40+yG3GL8lLsQ13wZEzmtKTW1fW4AzSEBIUsh9+6QNO5HZNBUL7gfsk9I/Kms5sqJoUT
NiBOsNScEJZRH1fB8pX9/zTLevwWEbG+wss7gRs1dyZzNVrC1lq5OY408dWyjlNJ07WM/hiHr+Eg
aEzW2QzcP83a3ShCdkzmdUYNZ4qH3OA2TzIs2KRTC6wfJXnu99YwAOpT4PdUNLv1wZeibh4Wd9zy
QxmxaA5ccKnAzwEkbavovOGWjuNeyF0x11rpa6Ub8PfQ3yIpUuWmVKVLV4RO25MUBQl9mgQC5uuy
iss0AM0SKsvstrQ3UUwMVPrsjI5g277ST8Ozxg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 64864)
3zZRlj8jZIvn2/dmjmOajFzcvcqUhYKgdUfHNSjkkHxQGMj5vfEe9bYDyq0dPs0mgrB9vz2MW2W4
hd8kTQZ/0PgJyUV2aAN0n3+RpVi5Wy1ZCPLqHv2iXvpgSfQXVKob825Oy7cclbrnZKEql3YpuLs8
dVJV8/CjRsFZ0euAx5Re3ydD1xKZBWTPGuauxJWAHDkvsXtJgc72tayazlzYdyx0uX6conw6/iRm
R+cVsOoPcvaTRvzqnD9HfjplRehNbW0iIMjvgwRRCYlJLUkQ4rr/ZYQ/M/f7wNjhPkaM0zk89h7P
AT2P7QJhmuXuV72JZAPMln+g/RudCIw334GYsF9s07ilr8if9tvbAM1moQDmi05aWpkQwCwgzbKR
ZFYEnf6VUDjWgfzBzYi9KpJmiykFFRJryFiq93GVhhLecCbOkNWGryfWfnqmk10S72RgSh4LrN8/
9cqnaSXOFNbQNTkRLoP66McJhOZlpHHvhZx4RigC2K9Grz9X57VVX5JhtZVDUc+2aYXJnk5Rt5uq
G8x9sq1VW/4J+HQNGnrjm1KaTTG9qWRrELVB/1OmweBX2MlLFN+kMcXr+jqon7mqGTNRwRXutq6T
NN/EIezev4LzlY9SHvEexo5M4eEXl1iaJcHb1Cqil9bGb6PNVZXcxQQC7PlwuYlFKIPEZXYvEsZQ
ihiqaAHppdAb7fLOcmTZklmF+yf63Z75lF7u3st5NAUv/FlDdL7T5/yS5sUVB5Mdgkj/ND/jmEEl
KKvuuHNrFSmGoZlpynsAEkMnHBKlyVxhN0BZVXRafYR7LaBfRnM9lz86c+r9eNZdpZoYmi42QDBU
r1cLQ1KQU4neIHA8QZ1odLZwhB9MtllFzjlurMwFuoR4XY5rR0K2lfN1+33RXHOK4T73KSWiSCUF
628TySw+7pA7xQLa6F0Ra5CEcvy3F1IxDjTacx4m+WUae3g10lPx6H+vVjBiU3EcgW4I+ObVpKnj
JONLoNiB8OHqdtEeuKa+vc1Nv9NcRfaN57Qxg6ilsjiLXYqxMpQBgE3CW62OWwwZjhPY+zIdOmVW
dgCuZZ5HhRqdwaVAcmyfzZtNh2CrzMHWl5uK1EVHZ730Z47yIX/K9F9WGkOLWikjVLVdIo4l7K2K
Q8Cjjgq+A/HLeWU6Hwaci2/NR36VGkcBADODKw/aXgq9B+/CaA60AUZR1CVOZvMaZbawddtx6AYb
Lb7RbbBqZi8tfiYJJXpfg6ecx4Dmwl/ftzMuQA5LhQOqXXWpwCviviBis0/xqirSihyMXxrhRFbr
Pwl2pu+Fh2q23wp4kqwOD5SDGtK2TlgTBOFxzu00u9jGJL33HK04OBSPHSISCIGJQIczVXhNUuEx
Aelc5iH/YFrNhpNSKV7JBQR0gJRJVaUxZXqJ/nixResmEBC4dfDi6qYCj+zLL6nuQ90V48Z6QDDS
qzQw8x0zs8TIelvjqY/2JBqN6paGlWlxHDXqXTNrUhfOwvWUyb7L2p27UnqAKNXBKUuLHqK7Bq2A
omOTqShFS12/wuf/JNxhBOLCIYXc8FFaJKhsKv+wSQvvd0Cdp+rmeSftUNeUSKhf/6LZAOQ3MiCF
vopp8N2i5yWxvr6M8ZSYShGTDSM/RmkdpzTkx0OaOF+gNtGgpAJgSHoKBdZq+TPVxQnwf4uES2Cq
YlNaCcX3MkK/5vuma0L9Jyv5TeMFi4h2tBZOHiAEP/EAd5K7YqKpo6ZuTIC6VYY9x35uZ4aGrxwC
3AOXM45UtYZ9F+ZtIJ17rFg2Hjz937APJ9lppUoVhVAT7XezJhL7s021bQoIJNjVyf3TUD6ba/Gy
yy07mHLPJbDRiP0qRRpnIwFQ8RHV4gDivsh0t7zjpzdMBk2w3Au9TfF+20bqIddyJMUiVKpJGReF
98GYSeHUT45YyJKwUbH+eQMLOnFEBuK/2giHQpJlFd/+zgkbVeHZJiO2+YJYY29KLA9y6LDNTkrv
CrT7ncGLfCWOjHynMhrs8eOBO8TibxCVgwdA71WKzuK1azjYvA+3TsMSuVV7YlajBzUyVGPAITV1
NOfZ2u6w9BgVgVsByGtrXkZD+H7RJOG4KBZITP4AH6dyG9qZCxhO7RbrpV0l31tOkIa/iTRX4Hc3
gjQNLzAuuIkTeYCBWlFKy1y/gixs5nOD1hBQwCkf4j7Mcu9+LbzAYjFvuUGr4IHezRfKJHzmFzne
3yo+RfiRbDeyydSWTuQnAA26bI60XId15fhMB7c/eboX5g0SIGaydlrXC+s3xvNWesQ0Ub2UW1j4
tNIqoENnd66zkGeT8OJTnAznywbTm6AuHFmF86HoqmPwsNqIsYPsmNaYRPLdwj99gMXjwssWGx+2
Hy+N6TVSopDmX4j/hr9ZerdrF5UABQjgLhF2dKefEKOP/bTeaN6c00SMCx1wvzeoWoiieQm/SxaF
rnJvKpS/7DVpls5tQWTYqYbH/KfZuJaDb4p4qjtlvHKnKcPJo3ryfao6Nlhn0Uy7jA/YgDo5bmhC
mFf32EHUhMUehArzFap/0AimLG/n4VIeg9zNZS5Scndq2H5nVv0I2D7qkil2gLABYd0inG3XoCDR
BHImYj1RSppaxhX2goopSo6gQhfc0s4R5rUCA+D7xQ5+CBS7w6abC5R/yBZy2jH6RiIiT4p4O5If
IWXJyUFHD4B2vcIrk86Zqmwz2oxKYBj1kkRvsEtNRTk6femeQvM6qLmflttZLkoWJMgjvlzaX05g
DuuzHz6bpexY3ObLQfXLdG+P1d8sd4+wB5XLjbU5R+1MIakdRjoZIpYC6q3vGVa3vPkgW9/MI1ZS
xLDe0SsQde74V+oMbnomcdCFuAxsua8Pm1wPreZc8ItNXNnO7Z77mQjrei5x1glEbtPboKRThrl5
a8tihqSg2ztX1HkGHlauIxnXJ6n33TxTH2hZjakhJKrbO4t96MuC8pHZsx6ZE1eFzzpLrIQfS3M7
uK2DNKcSRADyB66N/UPi95noECY9cLpd7cbJxjuPVe8eN5INbw5xWuns3FEx49/EDkDi7AEUCb/t
LOQPv+T5K7S7l8liUVlNmX4ZZTb4gidE1w/UK7LfzG3KSwf+HkD5AGvPwO44dctivL4KfjMkvKq1
hqswGG10qsyfCryH6aDFZQtvN8pZVsOLiQwgX2Dp26zy+NgWkQS6/Y9Iq09EWCgIZ0DsGmEPzeFY
fVQwXC4AyqOaviGGydSQHi6L1joRSyXPCsg/d6KFe7/qHnvDGHNLwViF/rA6PVFB0gcgFU0dbmrp
ytOZ9wobnkDDEqlt8bqyH55pPtAEdP8I5GluY/pGphH2qF0WhXNdVZmXIaidBr3Qiuo+/F9JPMy/
1JdV08fwvP0eicoma2HYX8501IPvzNvKUgjlFZRbJVMfwy7RlFJud5PayeShCO0OBZ4bYJD6gu7s
NXO23oOWhyoMeRzvkfOt7lT1yXqVR7+fGDt6mblb9mqAFVKDouA8zUzDonFSLHUBO+HQYNNOHNll
HLKplSgtHf6NhHu9QWW03ykZOYw6LiInF31IoF1O9ScfJFQCVnY/nUw1EcqJzw6nPNwlC7DYyZ2+
vVIfSj7Lm2OsT/9nc2K5L3NQ4Efy3S7ukuV5jufAqQh+h76O6OgyJElYoxJ+CqsVlJ7Qjtz0Mdc6
KGIS/B+M4y93IULJ/1L14U/eA9p9F/FuwAphxw7vnz50MfUW/Ga+jUk20VydxlAG3J559ZiH6JdP
vcfRZz4WL6G8dsmM6m+abfhUILE9juw5F0W0clnqa98KSgOyJP1i+FBJiWLHxMuPufzLPJNJgeI5
PqYGb3enkt3ALHWel+8FuEXeos6t9v0x4sL8ckSN/J54+ZTHT7bPhCh90dnMEkZ5epqcOaevy0Zg
pHljKVf6VsM70R6KsiHsLsqtyU2SJuSpIZiwx42PpnUJDkOkiCzGLqMsta1WyUnYLERsImjX86rm
F2wvsce1NY2DnVc2+ltIjN5/2Si9BipO/OR3+t73v8ZeDNeO9S0T2Zo9u+El6xq3gIhZMBwHnqrv
BrYl5MSKyWfCGjaxtym7aWlsmdOz0Onb0sIFZflkWlYdvLyp3mjlI9+yjYNb2gRS4DnNeKns/LCE
glykovyOEXQE2iYiKsggYM516BoUJFEXZ641xyLMWO/CRdCv21NcrZeJjYZCwO5Yy3M6wDMVmKLk
KOr6GGJaqWbXzKimzXkC638paROdsRAYDXPxcwHMZw58brl2MHy9rBmkcyOFScM+20r85aqkVQgd
sBzoIDMh41hKoca3dlWPUcRoeapokgScjyceyiZ5xoomjmE9PIXl5v+eJyEXg4dag0E20KPnDli8
abJkQMZzyPj6G6/zNosNhnNLhAAAgj0SBFY7mMG1mpdzHH+nhGr6qJ84jVCVt8Dlsm+RadhD5rgN
bTy4k5u8KAmF7rG8mtTgG/4LziV3vjowpZRL3RgN6AbUEn5ucryxBiD5C/qRX36gKpeKaIZ83RlJ
zwo0OeIbjz2/e4ykSWsMj7khR6NFoZ8Xyu2z5HPPBKB+3VtjQwnpp6Z6PXgIkNozzo0IH+a8rfv/
DwR7pEyAcS3XFwF6+gAQnZCD6aztQpMyB0lMA1w7HMxrGa/qKxDBCsfuKS4tZXvnQm/tPRIMhT+m
ZkCE2nBdl7Qq5drNTimRY0XeLMFcbJSUNjqECcGq/1xidsrDDNA81QxUDnqqGh1ZwJGe4yv1/ytk
FnMKTuVhh1Miqnr17Mq48mDcvnmfALexxb65chnn5jK/My3Bhx2u/t4PfmSVkTJrxCzVL64dWtNl
X7hKuvL/Qb8ct03FO89rq+4GasKppZJyFlxf86mMel5Ohvi3/S7cpCAa0RaMjbLMoLltcO0/41ZH
p33LtRBkztDnKNEkYbMJBaIP9s+hFJE0PV/C57BxG9x/sFGzErya0/hvEHv7OdLoKMrQzR2RhFV8
lWeYfnVS+4aaUfEY40ZfwU93uGVvCPdj4uJZc2rrZdd2RyIYGf3SAnh8Ov8iiu0n30MNcOZHOyu8
E0c32fumktmBS3LkSMzDPcCWEnhHSRTtBfnsyV7xaZsCJrGo8mY11XCQAnMCq+kWMPyWyGFEqcQt
gsOLLrJgIrBE6cOW6ajGf1JqclMfIkjUif4oX63vBK5Ux4Lh0LYiiofJF4Ha0MxcbTS+1UJ0JBmT
fLNrrtpN8H85DKeE3XVVNjj+Kvjuxp98s0Syv1w7OzrZndnMByOGpOLuwlF/eIM2jGjddaFi+zV2
OhIZMezC3ieK8rDM8CvgOQjgCkXtszMAU6if2ERi9tKhPUVmKLYzsih0zSkMQgK5qOIah71LmXZi
9s7+HPncJshp08gtYZm1f19m2QtqRlzd6o/+c1rQMgCB6gWXiv9uxjiTuNLxR8TWppHxgFhl3WiP
jemLMu1PytaK+2F3iEEkusXOiaYJgGAkeJ/plvc74AYlAVOJYYvuSJDKUzVruKYx0CVvUPIusbWm
wXla1MQxOR6K7hQAImRUIKNVu17yx4oSRgy7zlW5qOBbGqloQ+Sv52SExQ92/Au+uogjQYV7rsFj
62cahTmT7AfyeMxMzaS/RMzpzZQTmxybACUuf5VN5mifmOjZ7GeMOi+doVr+MSowHaC3iY+d1T90
7oQtyV5PHdiOKqmtVrT5wO/9LGnqt+qOtE3a8Ex7Mmg3PEgKUCLfEplrlDatIafKNjuGgPGCsiDE
OTgGEAxwhWTuz3Q397gMV7WaETbdlXRQJz2486K/mPeBl4fGTiGEhXCW5gj5bZRtRqkkl+YiME74
8hr2Ep4envezLgcsoaSxux8xEHWWBQ5ybRlachBiF6oPl3vxu9iKpuJYyBrvfpmmbg7jnAous6NF
7TSV5Xw32uWFtmzNl+QIzJgr9WdsWMbB1eh9QKfQvIevyCHgmYW0rAr4vlUMTKzm2Omjz9+OmHBF
dUZrBpSWsNo+1IP5suL5Y0moO5zW3IqxxxRiq8CNQHk7nGlq+PgTB94At8xKUTNKn2imQEtrtgpd
ga2DDwL2af6COxcFrwN3G77EYz0hn/vXmoNL/R/un2Bkr3QWRBa/R5AklKV+dMTj4KuRAwXMV6GN
XStQRuE4h/QllMstJjXtnW7t+AxqgCZyIgjagH4AEePcTsx4D8lBwuThZe7JdSxkbqMMqYnNrEhh
BLoIqLFj++FUAnZw/4PNCEIGt54/lbkfCZVAUuxF3fr9NhtLJxc3HKcD6FDD3rY3NhaqWSpOjgVj
+Zp5VCNNKBLmpDHlBdr+aWaLoRU6yUC0xL+lpSEL5he3M4w0GHCNPhcX7hPTRhagj7A4jXp2yrwM
zmC3wdmBCpi7pkfwAoeAYTYe7NCLxOnqxameRDh/tkQ0vbWAjvQ7AP3IVxP8f0dckkE2l1s1Uxa7
FQ9kF+H+gAkk44OUr1i1unh8ZsYXIcs04khs/9o+85+VKPhcOAgR+lLXtl5b2QHaJHfeyYBBZZUg
YFbiRP7geOGa6JqhvQGjpY+ETByIi5PJqvWYuDhzFiT2SZYkg4kvjbT2joHVM+gA28bQPebAw0hI
GbfMGgWIGgPLsFrMCbetdbYKel93xbvnEiAoa+LNHjQIvAD/wYBmFFi9kfisRB2tPEi3iS3pATvf
ZE+/y6JaTw6QHq+frZ93ZggY//8t9ehKQsyNvVJwicDSQ8wWMnnne1I92Y4kFh9DCxUAzZ1tywrD
jBvvqtpj4ebTAglOqg/wCr5xS2uETsuS4CO19TabockqhBOozhEmSn2JMvj6PbZ+/ku8xro7AB8S
9oWn2y7dznRFavLYExOLCZvFCNGJG5BhW9pF5mw3ZC0vDszu3xHpaLNDn2sVnm67lr5dMtKRe2AO
7oyCm+eXoaF4tGuTBBKLsF3pYdxDeon4P1bOA+j2555rmqICc+orBq3tlhG5/iO618vYQzdegQVV
o1+o7Iswk+yXCAObSdTazK48wnWjXCEwhQvRrvhDamxp6PQnCvts934uNJ/h+8fALlNzqt2vLLB+
5D9pGYO961uw/GhfgO+GlZzAyzDj7qfh76hV+eAHNihBBeKQjUgKSLCJ9huaKMV3MgrImn307ELp
fPMSagXqxkQlRAeIEqaymacf3LnTg4MOZOzMhWMyMbdl/wCC0psNgYmgGec19LI8MQUtXUQE3rx9
fY2jCFI+2OI4L1Q8SH7kbEhGigpdnuw3eZ19n4pneD/EtPmj8IFm24L+yuMwNGUC98uiwVWed/Re
+VRgIcRprBofRDLNwhm1TaIkb0k+gg0S9KywqWbOqgImKqMY5Nl5H8CxrKhX5B07/jTg32xK3iA2
yPfU4CRKzwjb8QfWDX1GJQ9UECurpM5plWL2ysjWDoayFpEwpsPkF/ohmgp+41VmsFz6NOiDt/xM
zl3qFY1daeHktkcYCPTrtUCBf1lk7ombOE5QJxceyVjJVBbrXVFz/nE7dWAhx7ultruu/ZBhLzLv
FeqpMPpKYpSHc5xyqDI2thKcCkbEP5/CcVWf/NRkz6m4Rynbzkp+wUVhKD6DrlXu4wKXktR+BUXC
ivN8diafal65weVvTkWGJGVuWCIlLKGouJTNIyEuRzY4x0oshyrlJ/UZPtMBAgpjfnAdzl2YVMnT
8iho32764tAOpG4f1Sm/pY7G76spjTvGl6yFqmKe5jLvcYkB+IN49peepdQWqaVYh6a45yxSJXff
ItjAZ/SmG6QgxMtzcqPCIX7DXAn6JjLST1BzxAz3F0PwKZ4tkbaQhdWnuf84MTonQQNl5QHS4m/K
+EBmsEBJ/TqhY2s3OIN6I9P9/xDAV05LaYE8JrDwGGn2DAZzQKLZJgXxeWCndTUzuIG4p5YbNNY9
JwqoLnVuac+euf7eiefaUm4OS34H+gtMO/81gNizuXSsjR7kDctEo70eKS/5CYtElhvQVIblgNko
8gR3pTfvCsve6Mzu5qSwhGlF108X+mhmSEE5jyt+zx07iInZMT2D76oDkT7i6Jz1S2LZCu1XUFX8
oDLyPyh1I0RMC0kVPe6DHqpQ9U/ViHtltjvOTRVLML0H4pqti/h0BFqwOOtA/4acpi0fAuH5GAH3
+Tg8CT1RRi/5L4Te3pKhUqsfXk+5gbKk8GPb/BoDf1BRa+0r4xVUXr/E+p1C92kAcamgWUG7tT3Q
Zl7yOtP+uXok4NnOIi/6mp8O4JN/f7hK/UFMxu0LN6bbFwHWAmZVUP+i7bWxrkhDPeJztNrw5PZC
v2bGF37GbDNaW0wPE8UPQzQN4NzFQLxBZjYEzNjQfqM1KhiPuNXZtlRIWFg1Lh4ZvTa3MezP7WFI
NsFXIC+n1flkS/EVATAarflRsKk6TGtXGqlFQMJJEp+98Cjp6B7OnyBmWHU2U3gsw5CqHEgZr5D0
ZHIpAV6GQZrDyL37Os3ji1yiFbpr4RIG5+SIxUwUAcsbvmRsN2RmiW0U7gJGWfCQKMD28mPOI8SY
/f9A0Ewx2stOO40uW0dHaX56AnTPgCP2zHZ7F4msrH6EDxjW+U8EY1X1JMFMyvupqwulcS8tfvFC
Nmfn+KLqn4t8U4k4vPPWyudckqfqKdTF7YjLq4GrgTVJXonrK28ZFeZnbTDz7+wGXsyrN+rbAqR9
NcRA5MylVOc0xD0NntXC24bDT04ecWPQDK8JfswpOnnRRPEpgBOaEgsiY94uhgs+AqpcfFu1Jwde
3bQdC19Icmz8vVl8GBYz25U1fv6fNlF00aJM0Usu7IHh7aYI6APponq8oIjmpX1FAVAPSkjbigw/
8lpGRh95QpUgAnuhMby9ksjnpOADugwesGwQS4lH9qpkZ5GryPmX+W+p4pt7804H/CzFdhzVhtSN
DNEhaCIx47XPcClNjxruFK18S/p6eINU3f8nhl1r0ibajp2Gz/9yn/fAdMsvj5s/xVDU69ar8a7L
8iPdgh0lXONlVe/LOOpIQmKqEiUcwW1MvX8LoGi6LOv5DmnQ+e3+lhnw7ITCQ/slIT8zK3RvpZp/
Y4HgCbHAzstKPRi2ExT9+Z6RUNheZUcRrvoiP3BnsG8iVoVLxNhv4EOvXivXlqYUdyJVZHbaeLvJ
7FdkVAb1Kgpm5R2iJqOaqOmhw3RqMEd0ck/0X48FK7kwUtflzH3Hp5tjl09Z7Y3ssuMSj2JSC6Gr
XAyiWNVoXVxGAYqk/OWd8c2mxdxaCYR8UtGhEjOqss8R9UpMgP0M5zg8egj50pisU3vRm30bKIhE
6RUKFrX9fLhKDeEgLBjerUFKQaggR/cztQjCPmltw1mx0osDl+aaW2PJbPz5OXWQDACiarxYetub
shkS7r9f/CuOELJBIGnD9DS7FKLORUj/4bT2SlHqsNMF/V5qMWTpO5278PQdODaCT1BJBJnvk/9w
rytxUFC9jrtfQklVHKODbOZBdLjb+4ILiV50aPwvvK/a7dw9StxqO3X2BXVa+wr0lBX4Mhs62hIG
LAdN20XifKA0XJUGlU1DrPVjWhd+NINxtdCHZ7rzhkEIVreQyYSnZQiyrwADZ1QFi9yOhp2PfjlB
dEowAC+umptNKQMJsZtK5K4YVHquT6mfAg7IxoDdlj1gREoE4j12OAUTFLph6gnuKLfzVOfjIXNS
YY7KMDBdc2GInPvySlYuyNG4fhUOtoQiuPDDRd/UyCYPUs85qqwGyRT9RUTNG/wLruNAd5Vx9k33
3YzbshzjK8o3YTXq7yCCRTyTaBVGHiRct0gEe0jjvtFKrF3qNMydOMZ0TLeax1lUMeggWYoiImWU
XCU4CN95cooO0d7/IcVKQ2Ft4nXEG213+q9uzpNfAJNXKatXREGNC7KKRF5fatnh2DSPu+o/aGzZ
jutf7T0zu3O50JTeckrRnZXEmApSqw8WacYeo33vKNE3SkgY1dVOISjAGwxcJmnY5OF4+ou/6oP9
7jzDKLizelDKpMxjnjX0dAXeD0Y2DTKukQftEHG/mAECpsvS6HqSXKVmBVttGhg6Z5MF0hUF/ZPe
Yvuvbu0kezpzMCxLomj9D59peTcoiiUprUWN4xZ49m9RsN4Rcp+TwGll7qfv4tqBVXl2IjzGsZX6
Beu0QIaBF79f69HsKBpinR34/OEBngPLTEk4hklbtnt+jAD7mVJ9kCc1IYBW5TrMJYeKrDy2HXh5
V+ZRp7leZt7yDEfGr7sTazf4y7gAW2z+Mz/FJMBM2zehnZrWdpYCaWfUXcuQ5LyqvlTYhbYKdZV6
effdLJlqiqS9eq6/wpvMSO+VfduNQZ0aU4iYUBCXvgupjLM+g24nmzvzENuviftcLlCni8vbb3ea
+Z2YO8MPB/3mgTC1LpWBOwVKBVQELNU3StZAsdLAcTbNUthzIHKkX1BTr/aEM8BePHpsTdMBwrSe
8QJVrb7mGMcbMyuvKzSW5ghw6PFsJd10n1zyITTZ5BDhvEbiEYBDpCuhs/wyNIgIDMtvZ7uDw+sj
kl9IOt9q0gG3tPAafiijqSMGT+KJ7tWxcs6mgAkP5Xy1LxKYpRALMnUeZCdhyCEXaos4HbafySBX
6agWmmnW4bBo7Kqem319NLhHmL6DwS1b1/7oM2n1PvZvAl9e3dE/M2GOGuu9NPAoE/Mzs4Fh+FqU
pVBeffTMo32fyMx5M3g/UFAiWOvBzV8VJP9jE/HYl+O5vtDWvPcq/rmsNU4DFg8m2Acd1clpXQW6
t0/0xehOlbQfeid7RsoG89zndfE6WuxYe6cPBltF9Hh11PnToLGeY+hf2VAHVLPec73NnoWTPJj7
DSRY4k8DIi4xMniklizbMIUmpr3sJ+48D2tsBLJtF0LFH+AR09DU161gfyM/BOK3JF2mlWG/zsq4
2BJN8Gqia/EYrftlwpLYybse48XFaXGK5PYKM0qX3Ej372nTmXHdObgU+cnfkrG1bGc9wQ0f/83N
PuP/Zx8/qRx8wtl/5NwWOOr5N9OmqVos/96HDC86aftTeQDq7MH19L0Muww4CICnd5l0sP+Roiwv
xXgQReovCFXtaU5sTC7qaiYCdCbSog3vhXkc4GcICoE/EEDMMSADqPtYD2rG8fPvpdRVB5a30DNs
Dv8chbCTq6gAg/u8cgR3GPuZ0x3077if/8ksHimbjissoD3PgMnKROE/W5+CFsyRoYt5fTqaLEdS
V81LAj7FKnup4ylpDo64+5LmWDr4f0j0TnEWh1tFoyupekBeHGTNt6LkmGfO7nfpL+k7EGg+UbJB
3rPdE3Mp8KGmDQQFQUqUtsGVI7A6owCQ6+s0rjW16sMvxf7C8q36eDB7d576k/vztKq1ZRdcG0uw
aLm3luxTmeYXp7iOMvV3KV5fXx2oeDiXOT/hOqBFeBIY52NrmKGXkP+s0V0j2plzzn6JdsdjWp+V
U48r6nWR2Xz7dMYh+xGH9HBV9Q3mCJ4i76iYNUCZ2eBHGLnGyb5xNkx6KjzDZu6Zv+i6sD/MIs5H
V/cdmSOEvwhpNxcjYipeW8ocrouUAcIoNyvxipXgA399Dn7Gtu0C06KNmtMscWbRrsRWmcboAMIf
AEGz9A77vQ+5s9xwRo2a4OLu18eFcy4iZqcwIYfCM6REVbb8+xG3osxZdjvp8gLpxNf1DowqavN/
nrQl/87Jp1FiJwB1s77Ap1Gm/VwcOUDWsnYKyYSrHN1MqBgkP/pIUqSz09XfPzQrrPQIQUgYxXn5
OomsiztFlOlZP8KrPzmqNwJgNsrGZWlS/nByTY6qDDqUx6gPAwXK4evmTTt3wsKpvvNto9QaK2+T
FoTOOWaxH6V9y5b91q7lMB1B+at9THs7ihbYG1fTHpMlXvRyUpa4uQLBUSdrpActJWLGVy+JBW7h
30DKZLEA0Bmu3rRop4CC1VW64f7EPpLobKJFpw39+Jb+zRcjIMF7p64UVCTJfHtRpEhXuLRhGp29
OttnASAuWmTkLoPYOwU6HZ1bTGVTwxBBajZRo4m9Blw4voL/dHN8gzgC0BQ/9vOPjNyllVXK1Ijc
FvQzODZDlsJT5W5LvKy4JBXxeeWHBaXRUjndk4YnuuQ+cjasT5aGTpL3DHTFD1erw0d+mOpBRB/B
LkmlQFJUCjyej2TLBPox53vrxDAEdMaUh3SpVLiMoIw7hW2gyksaHLZr3TMKS30kcd+kaCrYoeeo
/auMyqq1i+G6MT1E13SEwszBUoouONPzL6YgOcHfbFRBXrULrmO+ZexZoCL6xu4oTvuZqnp9YsKf
xEbdE0phBWLGqxKBGEYLunvAzON8XMq1dRhzHpgrF53dCKmQxGETDEM9WnMIRH9/zXo+X0IgHMsY
jgnTeKZHY7Y3gzosL9R0He8BgADdJ8z/n7JtnygyMkFktrlDoREc0oKP/kjVv25r8UfC25WqX7Xj
gh+0bAOYHiJH+O9rDLtMHex2RWBl/Hbld1w1g9l2TuMO9nB/UgsPVAdvptLEnJ4SN+/oZEMe0l4n
NzXbnkw7XPlVVRaYQvIIJ+Gfe+eI0QCVUOarGwctfsopuJdLxnbmfrZPu45tldFl041QRAA/UAP4
EEFAA3AzdzcbluLUtzX9kAqbCdQ+aaC5aK3i3P08E7svpAvo63KDW1bL99o7CYZucrl9IP4FmIXK
CCQNOhmjTDpusizJNIgrwaX6xjloTyWeUY7FOB94NW6utjWi4TAABl5Q7r+istEnOyaG9zO25nV6
iTHBJRGXARiqdcZR6kJjAfUDwVNbVOp53lSSdvgP66/1FJz1nCU4lxbVqyiR74AOnSTXDgOmstsz
+aKhuKsqOiXn29cC5hQSyfqVORtaTmAWUqBmECvLMnz/RtSWX1eHeWxGQoG8XytcSt9kd4H7+S1t
6hy2sz3w+b8pBATdfGXq2LF4B1gueb4pMZWyGQC17QrR6yyehs8vi8dEJsGEngAWxzDAuINs5Baf
a2M1ma9BvvflwHCP5m87awxNcsWTIiH7SZncogWUg7xHBQLADaQSReEumzWDbe0cWr9n6kfgPSXf
v1KGziky3NxqW88dxoGYD60uFo9JEjZQBse0T0alSGGjiyJ0C2XYf4XLecgAWQLvqpIxAxVLP0HE
oF5XVmKCqA2MnlyAOY4PJghnTGjSxg+f2lrQByCN8SJXYp855orLOA81Xe2ueAArQuBH+W2kes4x
UTOQUproZnmavRSK+PCOl5HTUU7WTVAt+cPbB3dYCKiMh+iMe+0ytK0tXfNie7NdUHJym991S8P5
4qUoEm47X9DWGFULOXfU0AktdkxrrzNJDRjlN9uHYz2boPC53QskcZZJDQQfMDo8rAh+fndW60HN
+wT3Dr66+YDLzv00UwIZh+UvCJg+LQT8c09cis3+Ytuz59Crv23N9w1pBcH0EEkDijnGsDytmii+
wuKe1Z4nUFBFnNIQRWPAbm/44Gi1owoKYruDS/jBOCSGn62sxPcneYbGeWSl6s9ZmeQB2HNtQo23
N3pwsSeHz16qV4syUKdLgWG0/aWPRp9ulwPC6LhqlOWaBEj3lgB4oS347JMETHGGE3ix6gOHtGlm
D+X36U6Ra04L0qf5Y3Lzm3seRu2BCkwQ78Qv3lFWUKxFtZDF1V3Fn5qOAzxFFaGSKNfD+4a/zzEM
ez5BatCQ/he4jvF5Y/BtpJo/YbMq9903eQ9n7U82aXbClZCVSNWm7vuzEpmoMVDf02H4WLDjyPfx
yy+5SWUnummL8BsGtNh9i+gqMNHlZvVgUN1XzwwwNL//2K7z6zouu6Q+QP/15bfrmahKkHHmcQnO
CJCX9H5Bwb886uGIdN4EnE7VF7XuXJdYCQMJnGzBrwe7Vo+AAaUyByCrveOy3xM7jEzXKCuWP40M
fZWKKG+rkcrPFT5cZZXH+x0Ja+Ok9v2O+q14/Mldp7Cac1k73g8YISIYUOWHc0R1ozJYrUWdg0n2
fBcORGb1I7WFHu2xit+9+Xm1ovOW6H1oB1yNbVtBSGRy7PuwEv7sya+Lb5jn/SUqXUgeMa1ef564
kwXcOuELRNw2bPmtuBNQGOSUMPW392QkhR5ybEcDYVP4ay6SE/U+EMhi36YX3sBkrTlFbmrh7HxR
54Gu7qMrhCASxwRwAnf9/uwu1YofL6W6V/UthRyJQTMWLceRJUspqcL3zLVnGumVAD34qqAmns8t
R80WJfvX01Pa6F9s6XrmmecZLsTqCuYj0wgSeqbJTOik445p771lXEOn5US1aoQiUa5yDw2ToO5D
hKQ81bKxjWITVHqiIlSRF7fXfdmwAIEV8C0IOkQZ85lbR3+vBf7nIUceiHafn6DCKnz/Wl6QWg0o
lF4T98VmpJ4/YsFbcf8WTQeX9x4g0RJI7E1MiJiiMLXOHavox3Eic1MHvYYCwFg1H0bl3Td6C/3L
oAHux5qhQRdKPWkiEX/C+IpjihaR1MQJ9gKNYGSFmtHDIZueUakPoKTgM5g7g5Ose9G1AO/KdzW1
32mNZ7E9KXbyVY60uc1+O5sDwq+86y+WjaVgxSX1jpLZRkcA3CVov15R2Y0lbuHlHG0g5eJWp5Nt
vc7hrLp9rp2+3HeFoAupeGzVLvzoVLpr2bEBMnQYykGe+0dpPzOHScFdy/y0Ip1jx6cqdQikVQBD
AVpCvCIv1eq7W3kb2udvlK9JCgkfyKXC6puLbdrMvK62hGpN/r09wgGrUqEQuYgosuBj/ACiczWf
h912aQtZJVwds459FI5j87BCKdINAiGbL/0f00lY2EUwbwjpf9Ua9pg1I9Nd4c7Twxvv8PWczWgr
oxcNVrSfvfsvwPARMqjeTDBmnPwfzxzkrL4BraElSDWH+IIF3x7gaOldynwWZNGXN7qlf063OI/O
i7MqIG98Q/eqgvbHYbr/TNYcnzfZam+OKcMhZn4qHYgZ2Ik6SpisHIjrF1YBUPXPClzXteBJXlWj
BwP8Oiam9Hu9frZrUMEC/iU/0CAZkz0YokK/rmNIJdNgHza2JJpLQcfX9ZS7sO3xF8CVhR3Vp9zO
aNaS8AvDz/l1XJCpDbRVSJ84T/Yykrdy5pG4+cOCV5I+DksDmA33PidN46yuzfwQWyyJajXtTCSG
d/1L2uXwZz4fFFvb/KaOSIFG8K9XLiPGFTb/qHo9/mrsHy4KRT5vXdURFpSba4jw96rVMY0A6y9K
NRezUG5bkyKRI6lYFNjcepFsPwq3i3QD4TjTDF3N+QpFAUXqmqlmDx1vZh2uETxPstwAWvyZGYUP
+4VKh/qW9ec0+T1Ie68Nw+blDBQJ2IsVnH1y1ju1+To8FL3DrjJCuxr511WfMY3YCitlgcxHnJAz
hxjzmukjpIUktvoNXGwIiGhUb7xKO5g0CnEv4N6Y/wAxdiQHqtoJJ909am9JnQ7aoHcWYtPj8Dbi
Ele4Zoxn83cKGPaASvtN4su05inR/wRVtoebeDpocDgsQT8TUxygGaJtbuytXdTe3zef/4NCynke
P+96q1Ie68ILdZv6xXIDvHu1pJ225Eycn4K2pPyAJrdnukKI5kTL9ISOo3XNifS1HND39mVAs4QD
q3F2kgLnTYFY0ORK9lbppzUKUK2GnDzhq2jZR+W2rDH4dXPMSmi1ybhLre36jKqHgt2RbAEp9rzl
kwHjoRHz4TgEymrQGUSZKTqd/oMgvWIzllg6f9cihIBGbt/OWLfJ+S8sLU9v1/l87ofWxo5dwIeJ
L1QOdhtond7wXkgWfPFhQYMI2wwzwltx2eYMTryL2sMmEqlJbNC28NyRfvjivMVPJzaqY3iFnC3J
ibVDrqoktnvCGhEcX9ziNplJ+Fguk0i4KJ5G7m1UmFDVPRKtq4WAXR95JmZoavOaGabWZhEyEbih
+/xZoF58/seZDZbKS367P5ZVMnuHHvMWqKsk8m8bDovkdidL1yexJV1QAnlJDC+v0QmyQyD5llEB
XKwTNYu+AbgUT2uqG8VUTkjFUA4HWrApdHOXmK1ifQySksdr6UQIOaPBLXNohjleHZksUcIJPIlP
dggc3tcwbDVLqbZrV609d79X3gOqAygU82bxHeP3fjbHxql4CymesNXetOYEhviv+e7fmX95e5Lg
m92LcNOMNXPfnDeoOmhT/MrnZJoVzEjtrmr9cT49ufKjzHbEl/Z1kl24spBQ3bU5O3D6ZbNZ2VIh
CgIaYXo82JdMojJxQqp3O/zZpKidA7gjOoIar4WyId1qhRxYUbvpZQe2IZuOZ/2oEAGMQas4JBFo
lX6Yjmk7QPtjemSx7P+nbhbR6OYxUq1xYqECwwy82l4IQWqAb4yU1nr5QTsYzJ/lG0fDOg1vqlT1
/vWVy+H4gID7owmjL6JJkYOoKtP1Tox8y79jKla5lSuC29PWLU3R9Pl2dCMSSstLykDzgItm07z0
U/5hMmpqGw0I3Jh3z/FXL9FGkDHcxS3Q7vGdSMx4hkBUed9xxurABcrLmFAjetmhHrZu5H6ESZrR
ft44SeQVh9tDinAyRDDC2rnxPb+fV6focs7Q+LRczE5NlA0Iq5rTJ2g8kPvs1XaHTfmR3mp7uz3o
bTf2D+pLHWKXw5Kynj1ZI1iNOBnk7TEYz1OVFPQFf+KFW63RhZFLt4uSvPbPopIVD7WW26UrOxpY
pbDoni3bc761OFN+BPIbeeGbGj+PvKW+5V0LM+Hayp0pA2gWZ7G4Wcb+c/ajRYJ+b7aBmk0bSlze
uCvajx1bywo5rO4i7HM2HGlnmTqiE4gomw5W5Gk+XF02f/7OwYU3pngs3SWI+Q7R06y8GvLlfqOF
QI8u3ft1qKOz1+oHKz5wRxonbLS5HL0DyVAsxtdfYwGbHmkC7fMkoeYUus1poxfk+Vp+7GqROg+9
nAThID1GEmdesC2PWfe52A+G3AHgQX1Wmvu6+YE5uSVIUZZ1qj3doHUU1PjljJXK+cQUPtiN4VwZ
SfAx/LJPjs+tkwgQpOuhG3uzCy7DH5X72HGBNo7LJVePjFZ+EAYnv0ojVlkUubGsQmChVdgd0/Ub
Cx/RyEdN0qep0x/lbyTsl4bmw+dqqRmJnHWWMfKdboyu3XcpnQjd47Kz7BZXUm0xE8tIeCM+xKLT
t1dSneNE+udGG5GyhcScHkewF585Drf70kzTRBfPItH0st7pzXeBceD3jqsKYtr4BXSNOdBnxmd9
2BKehItyTlFrCxWWQ+TW45QZ7SrU8eHgWeKjEpPzzp67ANMz2OZZOu7vBGiVVLPCcXUCvr+uY+GB
wWx2++Hs5m4L6m9Z9fNxozRB7Cl6Ho2iLMPstuWeXYjEd2ZMXk5zZVyxPZl1ntB3DVivK/DOce8o
zurJPJZlDjKxcm0n8NFN6sOYL2btfLyb88Te9BsO+aTX9CIsWphUYBuf3WcB0VuobWiu/unM0+au
t+zXQPAqNB0o5Lrw+dIStu1/a67KXZEguNw6+MgWeNir1/kOgm+w+toRt9xnO8rnuiunPbB2SU4b
k5814nR4FZfoBAIIdDKmtWP40qU0nzQkAvtELFCWKy8A/W0eqzT9RXJWVqUFn+CFSUdYkS7SJeRS
jwxc8BqVjfRQOX8Sxn8HBkDbYwr527nva1pG8DZ00den8m97wBixCO8DeRasO1V4zueS4TZExR5G
fIAqzhgIHbUZjINDL13zNm4vpJUI5oyrFJb7APtAu7mGF74BDj6KMdC89FFRzJ1B+cGOa+eEOMUn
CO+ngj1/POCMmiR+Xse6DWO9v+rtRj5injdLCmhErjYgxZQIo/7PkNEAb0FHn51EnqU+AhOTqBF6
Owbo6w8shoYqqNeiB1rOAmkCZbgmNUshHffOi7Wa2zHE/CeCgcPo1SUpvN/OXNnBNHb1VCFalmzw
6DiyLtaTIydX/qszRvlgXk2NAH470YXsvwBb1YskIyMcnHsTxYhAEQJ+eNC1eXCgmOk8ThSt/++Z
AmzHcuZnJMdBuN9SjUmmCTFXDSHw/eQz3HAlf3OVLe9F8pLGiucYLF8BNz7/V2QlIrA3QG17iKTg
Vlu60WrD0hmFJd12WlIMV0eBrR0ta9dXE3OkSUCIxba8YYq10B86tNcQHUEv6brpqLVY5ivg0cRh
UUciHGJhi6Af0z1XlzWWpAlIDaqp7A6duce8pQ14Zp0vMIecPnpvO+ol0xqx5NXuNhx8MS8yhOmN
QSXuQeibVGnChOq18RMQa4QC3pNwIa7EOY3WH8Wwqlb+92tb1VEEpjqzRiA/+Xj7qh6xK53A1VWa
6GVgFosP9pi3dxXH3cEK61Wl1W0DqmdezoZFD23uNQsFLEONzwxJAp3xdlPauPri918+zjAnbJv2
KM2tUkSJeARMZnFRKZDonk9e229ONOVzeYDsNVY2ngG8AIgflA7BKJ5ZsReYh8rZ+HU1t/mRrH6N
v5ZvyZC4Meoe4sQxU2DOgLNcBUri3Z01LUiIqXzm3GrPmYVcbOj8V8MqUc8XwpzdHjiGrmk06J0W
srzKxcXPwAzaHiGr2+y5oUD6rNeqPYgoRvmWS7f9UN/4P4GQBGfqpn+Ybk10MizP/2XNKrl0KMHx
R/Gf8+k3F4wS8nKstYcPCW7fhGqN/ObkNxLN3lVsEd/yrXP4M1iuWEQQgz0tAQ7u7H2Gf4tPJ4HE
5mTHCjIat4vqjoly1yQOe5HWIuGM3orCJVNBNT49GeHXb3TsfxNvuloxV7xgTquZ41nCG5/P7u4t
Qt4nKqW//t5S1gi/c7Wl1HdiXbNJ+XSUOk5Ln+m6RUnMwi7XkhuYBGJjfFp4COxZvK0LogE6WkPb
PYQkqnqQODYEfCFgeLpMYXIezXMON8nkNKseB9DkaWn4X7MM70fWJDTzMpJFV5XUsJEQBK3sKTFl
3w7U8o6+S1l/XwAtIRdWDQNvWbRaFD8WGGBUbi+eTzDAb8E6FeIAadBe+TS1jgBvIgwsRrWiA1T9
7EDfc0GvVOarElecHbOPI9U4e/XXZoJAsdvVAPHjgC4iTOh2pNdG7rIF263Xg/m2Z02v5IYVTLyv
RFwfJ+wSAskRb5KgwDLUIxyBfbSv1O5q/WPTdLGSoaZcAaejqsZMZrqqj23zjKWbEBTzcmZGKa4L
DrB8JAgnvGIFMZmRwPtNB+VQ0uJl4CQu0h1S6q4IcnPaosIOgYKO5Y3uq/WEAE1EmWgwtpAU5rAO
MdanWS3OBGOZM3dTbThitTqg8+DjXIKHnPLVPnM5rWVqC8398V2OSmbkJ0M9wFrTF4trA4x/sBDI
ZI5edK+TG/Kk9iLF9V4WzGHuVs6fn/qwxf8J5Ebvf6IE0VP3+c4zSdSfs6mJyDQaeljQX8HrfCLZ
fQa4L9REsDCCGAGpYhcm7EVsG7cZQc4LoFgq/ZWXU5fOLbdbhM3Kg2GE/uFS+bEoGxvjyGRqPOhk
w3D4R9lLLNi3+hqRaMG3JB2WmMT958p0J+wk4sgnq3+086yytHO7vy2Dz64dmnpKaGAvuW13xQ6f
K2OvL2+rOkQmBDWhrC4+E2Lkq4WZfcEmN9cI1oy26oF06nw6uqxLgtsfOnoHCaX1VcmvmwFsUiWD
5fj33B6zReZJJ/CBKIC0HMSn2N0CwollG3ighC7hc/KXQBUuidnoq/NlOVsld8utwqt/PdpWlw7n
bPJiEBZrcIOUbY2Jm5Qts5Grv+IBERZLRzrGes1kJ7g4SYVDJQ2akTvkk8AKuXZ14RKw9ZRXPb0k
/QD0kdW1BCOPbBkjeD6TBluwja1rqlo8ixmesENVy3PjT15DJY+ZrCgABz+YwD1kIUxZmliQjt+5
md77T4ExJtAqPUTJPsDYdNkCZQm1N7rYCbCs+SlE54lmnXOwOgFrC3s3frDr5EzrCU5Kfu7I8PTl
yCfJxxnRbOkadjopCaPb5rDIBiXQ7abHngfCguGnhEFNJoIfN1Vm+ZObRWdLHrUgZ0IbCZa/i8Kq
e2NJGNPi2gDgZ2xQ6UYtCqwrWQtljTtmhrn/6xJbMJdntEIT0h7QNmQZLgwitGqzBN36NXM0ewS3
1bFxpdwYbqQK38y+Y1tx+nrpEiUz6In42/uI2wwSwuVZX2ae5zX/VjeOyho1q7WhuoIhCv78Rys+
p5iYC9FsCr+jLjD6fCBMg1P2Cq4KI3Yx8JI+1faRFYsWC63pB2Jt6MP21TKN9QvIJObwr7MUVdt4
QZaU0id6klBMivrJdip0mwvlbZERKIUSR55erlshtB0H5tF9jDh0c7LVcmhmI0NM/daAUO6Aknxf
LJWrZLWL4K+UhkpR0FkLLH90hb2x+ESvv9gySaoItKqDvJQBJJDzA5Ia7raab05N9HflvumQOTzQ
QdfR72ELFedAhKVEt0cJ+NNw1vbSUdtRMmOGNnCybM6hhEZOvFEUNnIhKxGpEuz5KmkdJDAaIkVQ
NWZ22TIUNrHZCMxdhTZYHQj04n7npWEm8Uyf3PfV9OyXhn8gyV9xMbOSp7xJmweKc2WVMUM0HO4/
DPZwPDVeYB1jMhvJCnO07I/FPBQhz7AK+KOIy7xQCopK5d9ix6YovMhacVmHu2jRnBKWbv93WZFy
JPXnYX170Fv5VuRTErFHabxWq5ArtXmQSNdxiYoCOJFswx6+Vw3M8n9c8j11ycMZZ3hgGKOrqJ0c
iFaEeUTd3CghyKa/KGO0/dw6L2d0iaJTDYPkiR17GgZFOPeJuXvFYGZlpqphsqW6gYgcBApBv+DR
JzuxrGBGUm1KSGw3kLrBO1qfuwfza1pmLErFj3cKR3xE7lB/FGjlOor3/oX7iAHDYEWzFSg4l6zZ
F+g/fZgjWMr3QRx67tfTXMYjA/HDfjk0BNCHQIvEeDP0jT6E35UNx079B+5QGYlE7/g/smcAI4vz
YQXKHYkEb+cbCEQjsygD5L+kuBUyMCbTQNEHj69AtYUTc6p7qZqNjVlM6+7M5E9ij2cG3J5v/Is1
la5Pimet2KRNm155Fs4mHC7E86lDXU3k+WzjEfxodKUFpnaZghm8+r8EoVAlDP/uCws+iW7ZQWa4
Bow1JjgZHJv6I4zr3vFSj4912iovjaXHPzZT6mI4ULdbkMi1NumxalxCKfAnsKmjsCexPC2zB5oc
l7JxBDTOUFSS88d2CtOChLAXzBBVTSv2TtFSVoqgjiiWUTy349aieJrZDNhnDD/EkvgdSQRmeygK
gR5gbBDHmdVvZ6k6tm73qSd2gTxf/iq/mYi3B8EJYncX/+PX4WL/9ZX9Us+Gz2qllZcuwdK1xj6e
o2pEZ0AD9VvENg/J1icb12s5EMrLm0LER3jWmNM2Td/3j3M+JiFq7Uhk1qk9BXiAkdlUSop6VJbt
C2ALkunDygEFy82RyAXla8QiGLdAbhydf99jGb/Ic1dK1Y2+fwIdrlIaf7+JQXD59xOLd5R3ZDsi
y6ksJSyH4npzsf2ZtBOFGbZpVIzie5+eR044HSRc+dsSaOTTbsqW5A+ZX3Mc0jPMf96MnP0+Tw8i
SZqwIMDVNM/xbCEPD4OJ/9D26JpxkFVz7a1YxVdRLBDFacRsqvErWPQvwNeamam5MbGzXnncfun+
cRSP5jn5gWzzbcqmEKjUmgphEbFg3j25Yli26VM2L7mfLmN2L+P1eTvJVOsyPLX5PHFEqfeROwBi
zX4nlL38vMGOdp8xjtWteLZycqIJoYLfPrJxDdT3B8Nx7vRBjYfIx8Q65IQf8RuzoRdMcOxOMArq
5NC7hrToZ/SkvECpc1UzZvuyXnU6+oihm58lyrHa4aAQpIlOB81dO+086rDWC+aGrtyRdHwDN4Yo
8/lOxHTLAwwsWfhp+Ua7+6vVyzYvxtVE8T6Ap2baYZ9RSSCYlX81B97PY+D23iHno69bzbu8e7rk
nEOAJ5uKm2dDmbiGcG05s1OGHQPk3IgFE0C7lTmlDVGrIHyWE9tFz1x2ST9iT8Bv5IN6Dcr60foF
CLuc/gURDF4VYGEExH9YoSYCjfdGVfKecexbnJfOYTAaRbYgsloZWNoOrAnM4+ie+J4hybCT3VBO
xi6pRWj8RgUCUDHPL+oIRqFYJwvz4Ff4dMY5nziC9pVvdxqNULm7f6vluP+yPD7PuY0hMkdce0xT
anOsZLkjY1mjbLXgs2c9di87+nrDKjvuSqbXBY21SVnNC281faXJEyy7J3+q/ANzKtV/Ad6iCZ10
mGYn61oNn0/gn36xVbsMR3FPoqqp8LKc/nSnQLwRhIfhsUgjkPwi/PE8oXITRoADdyRzzs6BDPV6
Dygglx/wiztC/VAuPPBlHep1r6+tO7MUzO9vWVo4OJej6Cw8L2pM8jw3rn1QJhOANTNSvNSPZd+1
vWPKv+9a6F7i+FERzbm2M464PuVV77B14OAAo1XY3TXVwa9u9F+R04rFE/yF5VtF5ym18Q4uheTS
Zw9+Y5NxMB2AJUBJWA+PnkishNKMVbOG7DjfSdQAgCBHkTW5yiLBHrzrs2B9Kz+fckV2CKu4hnOg
zu80SJyChyshX7OEfoGlCU0J+LFViS7Ys9Y3IHJxKAJcf/7ZwJkfByBZINYwGMsm4LenodWVEUJd
i8lliIaju7KB3I1dGk1gKrwEnJoiK0X8BYFhWO5EXknGCZL24VqhKYrmIx9W+tmC6SMuiTqZ4Ak7
j6HKozJ7gC1rITJETmD6RRgdO8dMWzHog/Awft81Ycgq0doxvSx5XmvbV9LbRGpS5wsMstYl+kZb
b1oZ+bw+ZdZtMEcLKcXEIjrnb1Ua7nWKwuqnlDsEfwD67heCwLCSTKlktuKIJslhO3MkNJi6la0y
8SB01e4I/KZ2WldI+0R1O0OPk4cl8WAqCroof3kLq+HWUClkh4DTGT0chMuu0X3EemQD2DoT7kmU
yNj4VFnbJXfL7HC1PCN1MZ3HjU1Y7sugpsNmev6Hyd0LixLVgOh67JycCYU+E2geBsdR9AEq/9w3
jynHLicq+cvUoXlpcFoi1IxvqaFNg5JH6Qy5FWINVxqHcZciJ2Fn70ou6z3qac/KOFn5mL29HDfV
1Yz9Hlh3hm7ri4aqHxmVs34lgDP26GiUenx+G7lDMmOXdX1QNRlTM3BUo9Qrw5f2MmGeTkaZ97Yw
5um3ZDUDA8Ejh4qqTY8OQDjU6AoLmFtWVf1OzR4bniTENUVXRBLDPSUGRBH2iZGldmPoLt11kyI9
3asacoSvref/SO2Pf3vrA8bFPphwOjRTWkc4d8skklikxMd5MTlJqKJLDven17jiAVQQXSZxA5ji
Wx8He//9iAk4HZQhNVZA3ceDTUmRvrk8P1T1APGxJ6gEh+KCS+PiHC/9j+3RzEhrK7aW4OsD/gZ7
YKG4//QsWTWi2qHt5c3QZowzZ+bJG6FuMSKN88V3rFCHnjJoZv13g/4MHlVoOVVOeKYHlDuYlQiL
W0idaWfYJGzpykEl6xhmRf+29/lx0AvHFP9YDS/zkRL1Xnj75O0lZ6W+vllcWG2rEnGDZ4OEDvN0
PgzBSvFo7B/RsKVAOTKeJj6MSGLa8v3tUT2SD6AFk4qPfIIPqsjwg6ebz82K1jiJPUBnp3eUvbKJ
ID1zQJeVFyT0nr+7ufK1UpgjBRmh23Q4TAGY6OFHaa932IWQMmNE3lpOHExC0YvnOs9U23KJUBdF
16YkfrALbW92FawEYGu8K4imMyN6G8HoiaVodPLQhigLv6XdZxKLOTBZUaeXDf5UhITeneqQK+B8
+/VN+e+3JNKTyGCzvpy25/G0h9OqhHscJfzn7/kGuDqHgJirbWp3G1VamBuYVDoaxaVaZtiX2pK1
PCFbryY7RBij87pePd4SklP5x+1zK/ev1L3UlvEF25OFM5WMQjTIbTBgkERs5qAtIKuPjm1yJWVJ
GOTbUCobqdtgjhI8su7LrUY3FSGhR7EmnkABGUKpkNuC2dgdeIuCvB8O86kLCBxRRY7OrMaoXchI
1lFTmieFeie45SbwWBHJay+VwEzFsxM8EycLB+++iBkaNUdMYJVrY+NDLLsHNU0RsN0jYf/kvIBg
/1ECRkIb7iOAd0pM4aHuQ2mT2S1Mpb68pvFvC1BB7riUoQ5+O2qlGuaG+B+61YtH0YvHkkSgadTF
wDYSC7c40b5jg56OlGm0i3X8z3SdxoOXAEHh4w11I0cIrtZOOd8LDOeLW9Gxzi5k/zm1M690STao
Z9PK8b06BErotd8rH2EkMjRqSpPIcX2lu6ZuzvMsoW/IYQaYDgdQq/9PErf5a8PdHGMElBfTUfN8
8ifFo+hnDtF5Zc06cHAG+gN0amlVC4yA6qHGCqZHevSfxL8FCUHBbYvCJ6fYzHXwHbyCj6uIgNhT
KfVyql7dBKZBcW2mhRUEb/7F/7/y8VfbSN7v9ygf2rmshX7B71rKRxfUkPr97IUtVCr0LsY85B1M
B1yrfruDjCeCzgfu5Di7oWy3325Xk3PZ8704OAzj3ceffFRv8PP0J4wIpHjbyW3QxJAgW2omyQRp
ieCcVvj4jIenxXcc2cCIXhjQUFn+eyBo+xOCjdGAutqvey2BHhr3gsCgK4RTlAKUy2Kr7vfnGiJ/
zd/LeZlUK4sdPivBBE2S4y9hM8AWl3a6jmWxp+UNZE7jWwbyIbl5wm7aEvfZFVQgmlfKY6fbl1t5
6KcW9fzT12uQ7Zv30e1o2P4HIJTNaIF69BsXBoXjQa0lrygWqcY70IfNAGY3G198YqSARPE5Vb5I
wYBlRLrBrSsvTY3YTtAKyV/OPTyBuLxg7Y/C88+3ONT+/2N95cRIu+ryWTDZh4UK5Fk9g3q0J6L6
uc712xLMmAW1K9NRYCbVvmCEtym6CvkQY49eevRlmMsA3q1Sj3IgEL9Mbdj1L8AraI+tiWJ3U64f
FpXuclIfnfWP9rRQCka4YRsCjAWBdVaT80Aaj0Qi7uO0PHq95ZwMm3wwPpaqcUUMGsSv53zBuSry
+iJ88qgKdyrqgMulevmQl1p3fHJBfcTH8FwRVRDRCtrLEA6V7/BH7fgljlSElmxWne+1Ax3qfUs/
7ZdS4oD4Np5ceanFg9az4OZjIXq7RKnU4dwsswQvs8xNl7gwwAE1wlHIcEzWfE0XC5732EDlH12H
g7O17vyILAGSGRCOCRrWK+FEVuCmSKq90IbMSlUioKCkuJs+NRy9ZVd6TPSV15I7NeR87WfeVrab
k+S+Mh1hCgrr6Ag0bzcrr67ghHiXPVHUD4uS5cHl12IZo2lS7PF+KJW8RsXJaIlEnBIuZrRZCSRa
bOY/cWJZ7NW2w/TQgfpP3S0c9h/9Fvg7HfmP63/BF8Auiexa8vHd0MgInMy9gjBC9+tCDu85GFf+
3FPiuhNFskLk68TrPhyko76zddgNqINlPYzc0qIyuev5ASm3g1mqO3ZqY/+TFi15kIVLDgLO2UwL
buC3ou5VJxtAkrpFp5Hh5e+yQPOfmusE0WoKtH+HtzdmXrtrjVilVKcqROeq9olzEhKPsCPlGDxv
cjJx4M8eEwUtojuAub5QQ8VZsmxgJOmc6dkTxS1+4jtEjtPRjtjGPr6ohL1GO6Zg5ZLyvR+0uhWf
+tKIvUEPGTJkkDNaSoBt96rVMkPWTgcCh2SrvrEL3vpgyaNUM6o7aXhkayX+Av/6M6frenF2o63j
VOHCJ05fNBRPONuiUghJPOwiSLHmLjcUB2SOo3m9woH+SjiUe7DQ9Ka3h1MFbJm0vEErbO4c65vi
8T77P5yaQVlTRlz86TYMOudPTF3Zz2KwnGGpWLgByO3XFkVMja9SB8SeFzgszJhgRgvDCUDD839s
Qj+H5SARgXF61g7mzdD+G58SLliwMXmUm/qJkBmk9G/Qcm8bTdNuJKqXA5i93UMsQRpsyn8Y3TWa
DA5pVM/bqTQ/AAlyfrQdvgU8Dh+/3BmnUSPh0YE0maZKWRz27PStJ8KrkKcZDHjzg9uvbNaTD84q
TALBd+pMUfwt0Ofvz7gJce8fuXZf7ZRdgB1XMBpySOVdi/ITUSxLDixkdjmqw29OWYEswzVHsFsx
+lyTEeTypsVamXGkavtmVFPVL8fqlOZSJ2sWDWwfZ7GPzmapb0OPjt4OUFS9gs3TjhluHUcTJyua
+FZubUptvSEdTizLwN1x3DyadDJetOX6TZy+1MhjORC78qSsD0rp0ZSeiPk7gd1FAhhn6brInyfc
51uc4acsJeYpgmu8OlqZT6auJozBTs5ZQqYqVvlkY5tZgPFZZVwZVN5eCz3y0hRJ2YiMTQxUSY0t
p7vgDrXNfqmlIgGmnubCov5ySZTt4S48qh4O0UeSH02dTjKBhc3ZxazebM3lkgNuO/qCCYFQJ7Ef
rRB6W84bnPxHRTzl0V+y7xze9wYzVFM3ybkBzynMIh7FDp5/vHTQ1yCjg8kwpOp3R0YP90RyF5fC
s/FdYwNVAyzHhJ+Pll9UcJT9657GhS6QP9k5t7YXmJxED/wvqJOcgcV7XBwHg1z5sBftopGy1VCr
nqXLKLlfiDMwehXbPaDZAX49Yk55X+pRb209CNGNJyqZY1ruDFIpC3vYtB7RM6llrTTZES1DihBz
IZaeskJ/bzAG+iaC9K67zXWSMBbQo3MopykG9ZwNbkc6CDNm29/Jq/9smLQo2hSsCjHFxItq6zHg
KsccYDZsGu52eYQU9FF8Z+5R3LJ9UxDI0fx0XyeumADQXeW6VLyoYFppBrm8o9S481Xdw51bGyaR
fiZktn2IBcYtdLQf7P/667TZ/wJxEacurYiMDZqTwG1j83vqJfq2J/baLZJofeRPZMUdOpusiUDl
k2boeSRwo2+fH6hmr4f+CxMyto1TbfzAqDdzYeGanqEEdY3HtoeJ5fBH1jRzgp+I3X+ws9ytcnNO
2u1u46qR44fnOVmDh9hhTqer7dw4Efvyom9vVQoSpM7MdEv9NIzLKMcGFDTIzi5K8jZMqJwQ4cff
SYU2pzXJF+Pbl0EWArUh3lV7XyMl1VeQi2oA4J/rLbyXmXjZrYu5nHIepyIHN5/RAVrqQlkqEIHi
B8M0b+GpjZbrAJGoCw1D/cosO+bZFPzDXowk/8JqTLEUgM6+9Clz5f8VgAmmuVEkOeQVqwzfIjAF
A/6sMLudNW1J7GSPPig5SWFaUld7GLf/gdr3a9LEOOCLvxNE9fXkhGVc+EsWFtsNFMeRvq8F2L+R
HOth0zda8Np1EeZ1s/mc4GkZ9PwbQU5Mgs4epjSggoEf0SiuTnarL09m8MT4paouxJ3GfQDy8ied
Xfki1BKJox0nNAZ09vnB95NRA4f5K3WJmTAMJGRyRYoKXLKs6B2wvsE03hNrlcIAH1SfBDNgvMZX
WKkslF6/Yt4/nW5rhgVM/6lGr7TweUnmnp9Zn3UIGXCLF/3y5qe38SapureJQEMdWG+i07/S8yMT
SaV+vNjUTIhllbjPoWqaA0lnxig56jNLpx9VGvEc/mTTQT84jQMCSPkFID4Ts/zm3wWg5AbBB7iS
DJqRSM3rb5D7HmLn3MRWtqDidSc3WJL89gqBe5rP7JNdRnD2lkEj7HSo/Xja/kPjVIBefDTriH+M
GOadic4eZJqr3C2msEELFWP9mN0+FS06Nx1Fl32XEdpULY8gNwDxVaY+699q9qIJLg5fLGVxHTpQ
zA18dc3wNW5eERz3ZeavIm7TDJ/LBYRAtgbPB6xwdOIob3p9OoF9CNHPXDHQFdXR1HoD+lHFXh+8
f56TGrNX8ZAZIoWPGDzY8TEXMiCbTWvEq56zDLVAOk/mAwha0U5ZZy7b2xLxkSUGT3SOkiudLNz3
HjgvGcgedc0DnEtNeRYfxtexhwZhoG9uXIxHBQ3DdcYCVwfl6PT2SIXwxLQfFKwTRwdrlnQiWyzQ
xW9a+cDEEd/Dd2RrUdqRgoLSgq/Of6MZ8gbQInyFliH8kfqH8+kySmN53TqM91Zm/7xBwwWEPg8d
Ggwfno/Vkj4SmbIgI45mG12JlZTlc/fMdd3r80YRxyimcgf4ijxc9O2qDxu/2Ipu9QRHUqfNOu1v
B4QE2X5p1eAZ9NJze1ODgVzIIpY/2Ik4M7rL8kKuD4uA5QlVT4DbEey9h8ef2Hl5j3qhV8vtnQRo
ER7266REIBbZsk7nLVF+Cyx84AxBoZ2+fKRZeP03qQL7+TxLJA3IgSnl9Nte521rvmFR97ygFUWb
ifHUiNDAYw6hmtovJzY6Xaf79eNcUWo3ihXcThxPAQxCwSVFVOKHmIdziQRzY38qaq6i20Cn793A
lHWqVLgIgQsCZQde9oAVx30Rje+MpoAGE08BixZQ/fT130B2Ss/2+FvoDwI+Sjg2E8lI/osiYAAg
OC9V/iHirstoWOl4HXijpdwcjq/+nmV4tSKOgl4Pc6MWzycfgA+4o84xDJfcEtA5VIvNmXwpFvnR
wMYypS26EZKBktqYTofMtb4lQfZqxwxyNNyDc5rkXHvmmO+R9jh1f2wyNF4hd2ZhxUlPk6Kul26D
XqY+5Dc40c97pDGC0PxXqXxec8QZBvzPTeSlyg9T2DN45olT9hHNNTijIv5s3I7Vrl0Gcv/NbUIO
1yIlCZMiZqolFGsaU4oMCHUUQkAqw9tsjlN1X18IhWP+jk7M0vaYVw01/DYum+TpIcZtjJ31XGQE
EC7HORJ8sBl/cx1EQKMo925Xy3cUEnCJLyotyKYhlqjBCiqASDCH9sYNEAg+S1wafgVvJallkEHg
29jPt4AY5RAFoOiSbdGmqdUujHt6ypFfeN2OQSdVlbkp6bTZzERIYJi0NM5l0CzXuFvvGzQRKLRW
Y5/b0I4+tuZ6oX0TLDM+ma84eZbJz6hHfOmCGUM/ZqEl5Dd2iehsn4PqaDvzAuVTbrVCHLdHGWed
kjo5B5/EwWR7/Qt7OZHpFwY2ijPeCEEeo3C5+RaRL4DebZdqJBb6mjpXfYcxGlSkWAF7O7mObDB/
QGyR0uxBWKLJXvh0BkzqHE6gUNCzJvKGDOeARhlFWs8yi+DV1B6JsKsu1qGNhKHrxu4O3ZKu81/f
eAjcviiz8ZIVuSlwbOptm9dhZgwwyh4Syh8Lb4AvqFeENZZVN5xEXXJvhJbuvJ4V2j1xBfaolWXD
Pd+GxCmAFGmZM43szBfaGxcc9lGjnLs+fQpc1mYqkUqxJRMSLoITt8zwLnVS1NWEG+SgE5FiA5w6
zXOoP35KYv2FfkV6XX1Or2UAWLPQwKF17urr/r49+jfH0rJ8Rfe8Q6DAdjNa+WPCxNYhTFaKclpA
b+5hi2wYTqu9HIBKrS/v3sS3rGyYRmNjlJjEi4nurv0C/Z23AgnUNM0sN4I+2UsEaa5VsC0/+QuV
kYobvPKVKmGXJQhe3mmPOuuUMbba5N3aa7RU7P7irxgh1ZLLaI4iMns3C596WhPXxSYNIbIvZOuQ
vWWHS9KAiXhyKn3hNzhYUx1ac9v9SOLDst7/JXz84C++ZeWLLVuHL8l2Ka8IXBIlMLJmMfmtukGs
zIaRDgod2dLbDVDc+z9NjtDQYVBt/5bHyv5IMq/pFOCnwO3eBlDi/RO7whQRO2Moi78AsiC6it4a
FCJeijZ2bGrhTE5QYXQOUlaWLrrEv7syi3/MhM/aJrjS3lMhVX44CoT9e4B3m9Q4V2J04ICjmU2f
K9Rimmy5FU2oRdI9mcZHxzPasGKp5V1b6n2otQu3yKVn+FeBwWB8mdWAPDn/RAZ9PGzugfj16jeI
2s58QsaRdJJnZutxHJZFzXeEqexLZxbBrZbH2AeZT8Uz6JKE9QtoX5/BjtmNrU/8eKcXyam6y/RH
n++M26Ar/VEBKBpvx2VOz5yShsoIdWwK00R23mY3OdOdcsqH5XXE2kEJjOTbpJC6+uWJbkMNwXMB
tdTi/Rd2bSH+thKW4vUCN9ENPYavL/hgkDWGutHoS8EnsWW6lUEYU6hqlwkSn5D+Rp76AILDHpFE
uXIEvSjt3NebYTR36b4/PvetNGzLTdnUpyqHP6E27M7jn6lT2wKDQh3j2cTEhE6vsTAnkwYnnnRd
mFJgWuwPZTsZsePNr3nOkH82BEhI//G4UgsCS0hueN5Si1wHKJR2Vcts5gsRO1urJ46ZFPmEG+EJ
OQmwbxZOepdM3dKcgS+GA88/hoL6sc2ooGQINtnXN0vANcHL0HAqE5+0j1kQVoxD6pQi3Q6Yi7LU
TyJ4j9YGvkXfK7jkSWHR3ZkZ1oP44CULxrMd9B6kP9lUS2aSZ+bOxMA0diJ7QKgTR3OCnvJv1E7l
AlXPHDjcWBzum5W2N3bnbCjSVxY+EsVpIHTWnQxEsPjlNNHcJHNVLyPmcZjjijYHcxyRsJw3rwRP
C62b8Jvi1uqib6Cy9RRAw9UBBWNUK17hCoMkA2/L/BOAwdNkq0ltRgznNDL6yAjUyWwLh1iGEoCS
NN7ywcrHvum37MrI4vNCpzUbULp1fwuR0n4NrQHmuvZvycGyV/OPhQw3dKeN86I9eDM/RvMnjYo4
R4O2BjkNCNo0P/RBg/Ttng5Yv4A2L7jd7gkbdDSHOjFRNHQlqT3rBDUnlLowIrktFgerYrc7VgoS
SI8tyFSYGIi+o+K9ehiivNBEwXp3qD/AlbdbIiDhswnqROg4YEFk7IkS5ss0tm+I4791oKtR1edc
Wj+CXy8S8iT82oFkorIGpt7aApxUUz5gNWpjZIVT8stWnidtxuxvCXewcCVRRdgRUCkANgSAcfDv
Spz41BZB6X8/LDcPQwN0emBfAr0+PV6SpIbRmPA07x04EP3pDLICNNiSOJFfWWjoTIl5s92Z1VSL
7EzO2djUw3o69Hdcwn67PUZIvapJNi03IVIqqqyOCQ2WcgfczrxkolbND2dkVE4soH81uaw+naAu
1oYNe3ltqCl2cbI/NXUr8V/S9d93OloSAgB+ECDmRRg7PiWMzF32IImBQKpGDN8yNqVUkp5r/yrW
JmZeVjB8ZOQEAAL7zuMLpb29zK6S8qQv2550yah1HKNla1rrR7gLVOfuX9NPPmFjLHHCNodtIMYC
bmglkk0jwiYY6Vn2FlDfgYe0MrCzCBwpmgMdmyc+Wy2XD7T8Y6o6eZnvkhCGX8+QF5Ml2nS7Zs6N
kSSs4LNijFnUeNnDyEgNc+yU0YxO91LC1k5oQW7p6x1cC67Hje3NQKEiQxtP/cIus4hcrJDjnWWy
DmWnhoIrz/in2di5vsPbK82mtnUshcyTNLsAABOWXZqVyTpiR+FJkrDFbISFh/TEE3Mx6WG21nMH
zZuxK02653VO2I20oxpOFDW9g0+nSrXI7u7OgHCs8QWWbE/+zSYO0WqonEqZJGmFtpKOsBo37wEU
cdkWw9noaC1eRLmRZxEjwZnw1J0amqPeRT0pHjWlJumWFC2dbAcKfWPwsHWOYzqJRQfXjNXJh7MK
ykjqmenqQRLddU8JHh4FBquXkwVk4Kj2b5HJsl21/FvW4UCKYrXDtE8usrkzYCFfD7ajoG6Q+4hH
YBxOf41txMQujRY6DMc3h3QIpibRZh4puftKqY0rIMHWJnonq1smYCXhMcx3KNk3wlxe/+CUDgX0
KqNMOmJSANs0Hu9lJR9HlqGW+Ux/4fLNHrnkJ2REbMTBH7OfcMKp+mx87+8IjHle+eilKCiTwUdF
DjczWq3cHvCSlwsKTuDc2/8pntwd5dxO4nzYSgabMQJqAQUhjQygf8wV+3oEcegFMZBxdMqsbr7t
8p7LPQt0QSR/IyGonW7F2vKTkL4KOv2PSPmK0idtXDDFtx1Av+LkcFUYJurm7N3e3Cd9TbvTNTqX
L/FJ1Gl0po1PjS5OHPVCb692p1s3VzuD8JubwS8lNbokXf6mCQx5zFX7uXNo67PKJKIcqU4/cYHE
+g7y09lxEvtcsKhOL+zcYkwgi68XgEfCUCxQql+TK2wsHMPxa6dmzFb3i74caLx3ijZHwVLFMHqW
TMEekue7HSa2FzTD4BT/N1BpvXHFFqyKJyFK7lxBmXM45/2Z9YnMl71QjmunEkYowY9zylv4ecum
ZtBZ9ydbSQpThOMABiL98YYqJxUlrFeEwmKCR+FKQpNstMqju9xrZdDgPlICGGX3YShTvYfnB1zr
EauGsP3VdUkIMBSVR2PdTj77Od+fjPSuLkXhSpLKlU4igZXrvbQ3CbEl0XCcQtT9NcAe6ukje0dJ
5pIMRmI8E/vIRpr/7ia3YEI7d8Lg11KuuAb3kx44MEQsizpv5AW9J8V60++F6fQspa0e9otVw1mj
kuuE+cVhlDxgllwC/4xpMFbommsLvRvPdM7x+Ey/IhS/1Opj6ge5+ZsSuar9/ttNH487cyVMzYVz
6z+tmORnNQvBbt10k3LM6+hztPNjCANmIIpGa0gE5lcbXPtCvJ150RbaXERUmWhnPPi1SoM868MS
ctE6TVvL6jy5Bedi2Bk59oPPjv0ucw9eTtEknMEMHEwEFownL1+RsUR4Pu1HO5oUVAo4pKwk9QMO
v/zzKlXjVW2eg9iXNrhbMCYQ4HEbsc5DMkxpViv5tmcqJlUBt31w3oBHcSbj0lNeDGRItZ+iPSng
2jTrimrHkFV4adc1487YxbpuLKFYG4lEF7FQlb7AqPbYOshS/yglkPUDUuPh/XdOialqQVIvRjJx
JBEa3AcEY7LXaY/EGaXqfbgRp2PGqtCK6mxfvl0F7156FD6F+CpRrxyN+8CNdvejsuAnqpACXNKA
ba0USSPf9PXGoIrWXsAHJxEP1PCHYGkN5Q4dX2RNAFtjh/faC4DigrDiii6A7mQyaLpYXsN8MVzv
Tg7y8ThBkGtRRCDyXk51LIJUFLiE/84VtyksnNTwOG7hmMR/HLb6pUUI8Kfb5T0aBAuYj0eHEo6T
y5ApHpSqEkgHxJ7lvJ7a+V/Z0C+jC4X/4owFmtlWQUQnUP6yIBGoD30s4DgDcbq52n1035yxBiZl
1AbiQeU5ilydVuuUFHRikxO/yWuqj7Z26VRBIr9CbU2xPklPn/hNABJp7HL98G5vmDCfq1kRVaYZ
LCgjF5oOxep3wvMts0tdrM8F1d+bFcY5wsomYeAEgqCpQCstsN2NBt5DfIJEUTEa/e34BPI/ptMv
HPjQCD02kQTgXzehdX1kpajBiuGVjOCkwgFhhPAGhCMEAsgS6qMfZCjmjrvTAY5vBnL5xGvNlsHi
gygOpIuWfn6/nnj8LuliTKwh33I9mGSTqAod5sCvmnSFVuqKtTSZBgq+DcQrV7HZFjLqIo2aa+Ar
eUu7S3kS7fzp9nIihD/sk81GQ2EcRD9U+b5aeIVLL63Zd/yVhgaiwI1hu85kXNMSpf7l0PXh31/U
vPl2t+I608CmQ0GsF9aM2VZ11pFHRrzNtt1IfjR5Oi5Iuwrbpx94Zyr9JY21wdLr+NaOpOeAdxMP
AOfdyJgo8/XBXVWV3hHo/Z4FDQz3nstVRR+stHvA+Ee8F+BDxPMxWFtlgxEZVSHIb8GwflqJeosD
4stQVS4tpWy/GIVaK6A94MgMxMfT9UStYx8aTFXEzXOHQUnNnA8vt+MBcRsgL8wOzl5qiqdr9f3D
uS032/hCaHsZV5BY5svK5EHmDaB0sXm1rQ7UAdHw0ydvg/eBT9N259FJGDcyKUUV/Tg6P0a4JTQQ
PlJFcH06zP1TTInZsZQFzjX/hkOk6oWlnvSdApDlPZZJx9+AeJ/qKfYUK+zdoXxPJ9Ywn/vwzWLd
8xTrpjBYEDZ6SxTSZliNmEMinY28LSUdrPZ7Zy+/IGq1E8lHmMT4vdOjbykQMDYfPILjoxH+9E+D
25sKp1kCsFlIxW4c2fSAnO0bwxwbYBVRvB/GWJRLdNQ383DcgVaVTKUiQVhBxUvCVqGWXYltTF/p
U/1uAjtWgkUQxKsKzmlKLnbCgOfimWeAQHlxe9ORbagSiT7FIgDJTfOSYxRr/6O94ZqFpObCj2fK
gZ7PWEm3XaL+16pxqkVS+PDbmZpwQhsaULOfYgGjdodWCcQus44LhXRZxoelMt+WWVftsKCuoDaz
E/FIwKit4AtF39eU2qr9xtRt+dpoiXYMRTicomCyMgUGzOlyUxZKkqa3G9r0WUBGdZgg5/OCoL4V
Blr0rQiLaijktRi5pAO7by7B2Ai0oFuRavEwyLrYrbCWgj+ONPbrsQDwqz19oL6i4w1XffZjybMe
tnuRActIubGunyBx3yocPnY6+E/6UZhppMuOgztEaZXxt4TYhiXW4sYioRvEe2FvHKcuc0pLIpEL
r6Adqkx4tpufPDeTnqj/EzXrR1NIA0cTyeGS0OH+uPy1x396JTx4p7MbgHSA/Nt1RofkOsk9YHtZ
GySv70ZcVY+PD6pKuRNCSXBQQqXoXAep8iADchnoUeLgER3xPqmOENWDq0K59NqZ8oRdBuwFFO0/
AyEn6IVpfD3u+MZTgZQx2pwMz6/k2yUNcY0tNj8VjUQDIqpwNZ/Rry9DCXjMtF4UfNoRnPjPw37e
sWt44kaAxuKXiF+61rFI9yTcCSu+JDIdjvY231EaqifjHlTqs/3W/DSKmPOZPJxzRNHtibSK9n+d
ouWkVpNNeJUR7Urd4u4ts2cirFIGAb8hc4Vse3ACN9F28aCfFP+tU6bfZG3HoqvI/qntY7vTCqWx
rA4kcywm3MhJMSGRr+ktiJnS4grMGIUuFXmBI7T5ggQT+/sLmRdLDE+wlysLbj9E7SEsoX9/Heqz
orqkNIaeXdmszSsU40NtFFZjb3sMkzhi7B1C8qS68M4ub3dZERZk4OzlmBz53VL7dyhtrV2VIS5Q
c5hFEP3eLAubNCzMyDDhDLexqAeFtdUK5dIdDPvByyLSDqykPzPDpZf7xtTj//46GfMRROrM6DnB
0fre95FVqAa6ReUh1nQNXBK8cTHyIQ1L762Q+BhMyA6a9D+mR3NF2lXPG1aa6gKxKnjfPSyj0zQX
Ds8j/rmm/hsId7Lpr9jEEQFNg+XW0KM6Rgy+EZbfCsl6YliafEfO+sYIbmce0HOm7JE0Xkq0SuNk
bn3+RJ2puYA4D1gzBbz+V8QJ7DFhY5OrAg1Esg5ujyC8g4k0v1I53igMYD62P1/bON0npJ3pvlHP
CKydFoxB7OAoaU5Mk95Cg8BmXEh7zfuZMawNqVvC52E8vkcVAto5qVGpO7hI/p+LPMkAiYrBW2up
Cn0OBiYaWKxHgAimrm1TnkSl3A9gOaaobox4lGpXGeZylcmmXhX8f/6wriNddLTI+vqdEvoOSwbb
abpkYMbMFgCDNCFookArUAOjJtQqgQMOcKalP5Ne04oB9UY7mAbL5E/aAWzAqhnI0KqTJjeM//37
WsZNYWEKSNr998wLUoz++RXUY3UZyRU0Szg/Z63ZauJIxG6zBGE7YRzhN4NHGPp3AXHauOBItMG5
0X/jrkmRQj3JAFImcnBi3a9cR81TLZdcKDWpSJe2FUsD0cJ2sHzixKcbOvvykpxPnZDZdtV5dYhd
FHeHdtK42ewbCx3XBq3fakn8twKuWE/asDUwlTJOLhGO0oZCQXe87ajrkw3K0FucS5Y4Z7rzGMWP
upEwGAIJ8iwr7ieslZxw0Ca4hvFM+0/l8Hzat7+NelQakLU1czl1xro8gfygHGcTqa4fGOD5WB4Z
hWUEd8ueHteQhi3hmeIQmT7xi4Vxz63iTuB7FoD6DIPNN9qdKk5WwLBNPzrOcvWOseIKc5DQ18r2
Fb5FTg2yxy9apiftp6sQOK28M5Nik5sSpN6DHbyCiRO/Vv+s/PKepS/ohWH0n2b8tjg3gxRfA4ir
7jCpGA28CRlEeP5/R6TvFOw4DiLu1vXfXsumdMrjsLS3QlUkxYxauDw74EV7weqZZA+4y3lzeWzo
5UXUEJjHeoV0O5onj89N/bcX8IEuFaUIgvqHJ/PWQuJdpfiahWFR3pBQ+rGDGwndtjCRQqeVinLH
6GRctGGDsvxD1MVLAtYJx6tw+39hnnhivhDBY5dPbmqiw7jMjXxyhllOj0FM/GHii+fW3UbIj3zC
OeeCCr4Cgm9ZpAizJmA3i4Ul5ceOlfYUBoKpvom6v3eJKWzc7AxEMgxfWcHUMbC3g1FF6MuosHfm
jvP6h+isCz9ggX2/HZwd8NmQBxAgQclekICTKlH7s/Hk1n7E6kkB3tRFOC49YtoCZQl0TouFcO2F
aXrhGkfm4z9fL26lSJVhnwldi5w4iXqDYXhyrTeiVyc/2gDd6EIiZBlUUaQpEpWVZoDsoGCvBcwv
73gEiahXaaUnzXwcwdJ/6Nfpn+5CeEkziSZOvp0qTsBWthkNRoeSbpSRSDYcfw5ZCzu9KO1F7wXv
H+SOgzZ/8oNtM4SQN6r0M6Ekb7ZJQWIgT+Laaz5D/pdDKQZoLZqorXlxsce2eT5xEeR6jVDoldBl
o3z8cAIEhCkP5cN+sarQvz784QlnqsvIijEYYUJ9sj3ck/Sw95DkXF6oCLN08fUbHM10dvwhcPOU
3Cro2E+EUj4RNiiTknP5+on/x9lxxK2uoQlOQFyTy0bzdEaYz6qinO13KIJpA5NtVGDO7m8SGmHr
SjD//wyKqPnGcWhw2BdytEbaUbLSU5uZOnhDgRubSsVkx0xCUMnPpbfwmcPJwBM9EpisCmD2fKPP
x2pOm+EEKJZaF9K9NJmuN1aumfKXl4+2S3xI3P+dwtTSgF+HkhHjPPFakA32yf6GMmlsHAcdvfLh
qRzFoq/VxQmi5iaHH/zQOmEbV7VVMTTQAjyF4skjWBQrw0AFdzydqlipS7TO9lGaVN4QqB67maFp
rfFmFTx9zPft9JBq7QnLY5uEFUieIsF8KJwbHrBxjECcuVu0TI6sajGgi1WK6Rk90q0ISRGOYg3V
47aBEazz1xbW7+F2y3V9+2vgYpVBg85esJUQHjOkdmA6StOWp4mR2QAdkIAH7eDVHuyMyjRnMyl2
RllzH3Re3iGaH3uxxNB6mJolw0GOgRpTTWUWaldofs67HHU0m+Sc35FR+PEiDIyww+Ke7dUAAAe5
rB/8eCv2Q4Sjnh2HosJpcNXBZcvfx1pQfSqSkHG8hMMVB3ZlTQMSpYT5mBVpMuK/JeroELywjUGD
FNCLSLfmstC4pzlRdmGct3qemna3z66MIpBlNnNVHXO8s6bH5FOmTu8Yu+8rA8fGNFNkfDB80ZZ2
E1b9ncURbVBSO7c4nrON9T23FSW3kK4A+IIbgOwWvKjWJvZOrEojyhTlOGQUiT6mYW3vymSNSyhZ
K35aMDYC55G3eAMT/wvj7vnUiKjqJMAWz1/NeQ0AfiOXI1XhU8Fo2ASYHARoBhBObEC0jVdA8Bao
ogcBeobXaCO0y9KWEIc9YQMX5BBzqw6TxkQYtQZ5e6VmURGuGzLjAVzlKzid6dj5aMk2ua4FChIM
3tIOGfN4K/mp5b7VxjkCsaLrZyauQDl0KQbiBq/l5mKMp0ffEbG3qu7eAhkoqAMyxeQodVxGkcnw
tJ5iRY5YMpxQPpIESIj1Fn6fH0+LyRmIevjjK2bhUObQTwQjzfXEvW1qm8WYpi57KZMM4pMsUN/V
PC0m7kPCgegNfMsnphU9b9CIs/vsgWXc1SuqJk8Asv21fYRIaL/d6xAFYPAdTX6TSffs9M7ySYLZ
bRNDDiE4YB4hUWLOPJNLRNYScWeFNb2Qaw5TyiOD4k2/gW0dn0UuFAly0sMxjjkab7oD/bGWNtxR
LDtwuxvRWK1eu3umlzS1ccYBgdk5JJDFiXES4rVwJ8zYrymW4qK5UaK+OhxjAIG5cZyeR62ehNSZ
e/TDksMxs+eZ6r1ODlsCchs/Zg4ekQ2mEAwDdf7hjrs+4/R8/nX1nGqT3LPU0KhatKQyjbX1sSX5
ATawqLRG360xZkNNGC4W8CpFjICMg1KD/rY/XY6PScBU/MskYZJFAuc1wSJfHphBpuiMnTfpJd5O
Uvmbv66ZxvSynuwRS8CkmNKCrcQyJ9tfyAu7ghfWU8hKHVZ9FDk794w/qolCOeFQpThmX4PzD7m/
qkP6HIjkh+6q0q1vxgcMWkxS1Q2AwYuWIVU9v/y5o+T2RrT1Lps/0NTJwXXGwu9o9n0dOxFstBqR
apUC99fXTOnamMbIpNbXoh9jIACFniYZnd2snJw0ZOReTTTaPAQLAwJE8LooR77xnL06G0D5bFIz
Nc2k0QoyqhmORJRuqm6i6DoJTFFAMDfouwV3NhW6DCjw2j6IZMsSFCLd41w1BxKaJJVEUcFBmX+T
E1pRvzljuqBAWpnVOIeJwQ7h6SkRbprYm2S6WMf+34k1rE6QL9i4JoKSztmqDjKWzHiNdUtDLchh
lCl53CL58J/BcDmY2F0tbgL39ZOw15X7w3VUO/vZhfAQjMSs05PzGoNTxVTu4MZNKrUBqMDKLeqt
b20FcIxSIThvGKCi1CLxAHAfAc5oJfdZsS3vhC4nWQ/U7qdd56VQYG4JPdKV+/2LVuSc6UfWe+rF
UgvpYgjebNcGR3OkQHjojjzYJJug1Q5JHm95MEFEW/2gi9q8U93I/z6vDkWkpR4/nW85N64vp+Sh
Qd3pT7OlphWkQoGru59BFLECYyPCi+bgPXfR2Pv+ptnldp9nzPRVK+6xzQql+saqXa1EmPwrerfY
LUsBMRQ/oDvV6oc30VY8sf6jkZ78yn17aYyjSiGNXHh+BHk1OLyZ2bStjCea8SSl/sJUSy4gwnK8
QkZtsmBS23STAuPllJeIPpQJrWXVnnqTiVWGXkDaeo23LkpSUM4Lo7BV4V57eVcUzcsb92AryS61
qqT/6iM5bzG87t/q3gf9Q2KDjkAIxhTMZr9I5WzhaJQC3gvUXH8Vg8GFXXbjARmq6XVo6d2xCX7m
tguNuP6B5cvAYxaETBQQtRe1ys3/Y8is2TKGRGLWvoeU6NPap/WabwZkAcmf20eRS3yiDp+fmXVZ
FOiqemXoqqjUsFETIwVTdBfY+1rWFIG9Ht0qv2RQj3QeL5IDMsRZsjywe633UcHSIGcd2DvI9d74
cd6UQQVoDD4H+LDKaVgeO0Nr2PpuF6uXajr2a27VnynDKdw2JhMbxKUl18LD0/Rkx+ALjVqPyICJ
N6k0HPTXdk/7YKJiSGT9houKo+9iDwBN65kyCDLg2/o1AFipnkVChN5YElGqOs/FvQxeO5H/hlMF
pwYWfLO4giQ2UwWn6jSutdSnCWb5j7Sbok6JvT+69jPk2wRZCgWnj+uuaqEGMarzhGkhd+Flts7h
Fk52EJOD1oemYYL+gZxNAM0lPpd/4lwYKy2gVr7/tkiHrYq2XUIrEWsj+RoRo99z3vU3JA8FZlyk
rQq8iMPdNcyTmorpidNa1kxM/vI3JZbZ/xt9bVnX8k5azLx0ekOY4s1WQ2W5SW4GVtPAIKFjeiXG
HDPlSgURDIlOqJi7RjNt43rTfXQVFah5QGs353O8fpP5tzJt7YF6JChGe3WW4APxS2uRW/6ReJIm
ciyTq2j93OlT1ZDefjQ5NNc2XDSkZZVVhXCH9QqFR9LPTzHWR2+c048eZJXhJpSwWKgdjgvwsu9e
EKrg58O3yOkBswPbzlMk6z001xyxN/cJbpt+lInw65JN+efndTxOL1ELCh/Z2Vo+unEe5z7cvOD0
tRXPuew0C4O6htINDSdidwChVxtW2p25vJtY3M7NbZAJ6mcfp2jhI7R3Mj62TLFjX7QoZUv2z0Om
kBQYSqLxZ/XMZwcpE99glFmi75IOMyRDD3mJAco+TTcLrAah+6O3EBxQBLy6rcTWtC8R7Uqt3yAs
MPNB3H3clhhkyfuT9Eg/wFT9qVDHFSsU6cJewW0CpCMmZPgMRN4Krp3P1Nd60XXSeFGjrJ5g2rnw
4vPzPI8TtQ3pqSPFey1GlH3Sd4W63juZin709J9YcCmfTFE/cW8yhoEfIUdjbu0jHvBbpk5ayAe/
H3ARcVSsvaE22TELjkBWPv854mQ8W0OBFZXl6L6yK0YIBemz8KxHiLRtAHVeVZJBy1hnZmZ4icRW
WidBIBQ9g2rtXbUpfqQzLbTQBsqT8n6RRkaM2A7S9K4Z5N3kfn0cHnbjJLsvD45F0eyyE6Hbrekg
ePqZzn0ehmJJrXT1XNVFR12fTuP0/kKWR7hAyONNoonGlMXaPKJbyldDHy80Oa/aQbkgPFZupqa9
3FfE6pbwTOpqhu/Wc55YYpUZ1vdZJ1VMq+oxl0I6rbsSumcB7Fh6BgbjgUIhTjH8mJf3L/4UXYJK
bWb4onSjXElzuL9k/++GJqmGOp+c++fBg+6FSkJADB68oLY3pYfootGLkBgPFPc5w1fb5uvMD19B
yqQUfFhKP3HnuapAe8M6mtTvVBHOuTsa45lqmcVddgp4PLo8B1QMqsgmn2HMzzQvPxgiPeKXaEeP
P9KljmyXmKUCl26UyBUHRGnawTcmS/7+9hvxSnxMB9I8EufKsi+SHZ08RGWB0Aikv0KPNQttw05A
INMeUeugtGYAsx2BO5DaxVxvhoPH+GrOpwxY96y4Xk8RDmXoz/3744GCNZXHkNxH9Yl37BgCl81C
31yoKtvrNvrrlTzxfbHVNGNvi4IedEU/esGU+gzJKbAxZnR6snIwHOX90MHAFL9soK/6a9r+KEca
n8lwFSQ51Y7CQyF5MMvhIramMfCtIL3r4mDVa5i9yCbS9P4fnqwVAF8qrq9R2EQLb9wcCHmBPg84
3SqXI6t69iCa6jOvcRt733rPRtbf3Z1WBJeLSZSL5TdpdUHhjvl4JQ5fKmEoTm+oqfgsmHNrourC
6BamJx1Do8lAFMAljjphrNoagLfKKeJ1HT4VbLhTpAwJKReYFe3kpiWMiCzJRjGOqJQg1LH6bbjl
ziIrjkFxanLm0NsnHWCUVjZy3ZUgqlazyc0NN3lwaW2WY1N8CEduPl5wm1OG7gIF9e7r9X6IW5nq
1jrU/cTY9yXb5S9r8h2FZRu+qQzoKNG98LaWxdyTXa6dV1dQVv9Q+fHwKkNbXz9i4ZDg/7hvzq/M
b5VUBDfesy3mz2tLEfzVMC/Iv+mvK1KgmlEd1vn6q89ap1OhMVmx7Qf7C2uAa07nmK+bZxCG8UxY
w4JL7PpuPhF7oFNngg2JADaWRGZM31/TMcYnc3ZHYoFAYEitOtoOTomizmCKmPs34QAXBQ5MIlqH
NQTzKGkBukvzg8umNEzKL6vMUvUJKPekImPnpZSJ35Bg61WuFdBZLQYBfsdwyO2zKosq2OUJ7mOI
biGuc2iBqzXe4dE+QH8vh2fOkHFbNVRE1cywdMeQOyAAnV/ETcJ7lzapZXmCZfllUodItKzouhQX
gYBxUlx8uWVS9nOYS334f9SQfYl6UAmn/4lSB4Zld/IAehuiKqefzvw04EXX1yoSsWWBv2Tfs37R
DJYb/EMuKmKE+GA/edKn46whvnSOIeg+L70uBbrBr3wxsZRaUF0/SsCUt5OMybAoOC63VQ+NGbOW
HViIfhUy66llj3kmFS07CbyNhn/BL24hz8IkeVfsrOx1UykPMxudsWkOrOtCwQt0gUTTyLtm0yUv
vsjWsupkj7LndepLfHSZNlszjUE9QRJacyvbILn38yydGBGnfI+3o1QvKIPLnhq8FmD1AnkGhxmg
jruAKtbER4wjtJp2xczzNt8q163ZpzCziJBYbxfhF4LjQO05yLPq3biVDzvYlXnqtHUqdWFtCAC6
HUPcS5g+LD2oo3iMb+qaeb8gVtVq8ptdpP/yBBbUx/vbbPwnhDWuNGYXlC+fsie74hsualimVWFa
7QO9mnnhoJ36EvL2sFhJztSYSEC1QAHbM6yudDx7SbuZVZrdb1rY9Ip8GrjKKcTJ+VZ7joJnXLnR
HG5wqv1p8jZskNHsZl0PgxMmQSX8vDig2Z7x2O3ysp/3bNgp+reoOweIW5t+5EdzXMXpTWXfym76
3T6G7WGalNhkrCg4bU9zZYrL0Aumgh08ZtZA95UJI/e4PInsVCvx9PxgAVK0EistlviBGLyQWQl+
D+4e00+nlsi3IU/Q0+SfaqMEvy8PP+SNPZUOpOhXYA92CzuBhsZV9XCp22t+xWZoy+X7G/7uu5Eo
PrJW/OjPqzbnMSD7/l5CZPR7TRTgRpyU5nxjwQOM8Bx4b/hHvSJineV+9V3ORvRMup6LJ8BPAYLy
/RUX/aclKe4b/VY5jXBZebTH5AJ6rQw+kc2J/Uae9XBEN56ndTPmjUuFknrP1BfZyELDeUJfX6Rf
Fl/F1HgINPGO0L+9OaKXewp2vSWTH4rwVhavGVTFBzjFTpMgwYCFM5L9fuJSakFztAvy+gWOPwKU
9H1cXr+DHfTz9SZYtEJ1mCuDcFkI6B8kOgQv822C7KqVbuV2H/oDSz2xgTmMPuWHkzvWDd4A/jHr
up0Xw2OX7Wrm5MFerMIbQtVIqYAA6826zdeqwaPrnswpGki3w8Az+rkbh0QVnK48UPChm3oVUCdC
nvAnrOm1r+ykM15Lve0vAnrID3fV9KCVKuRwMHFE+AlpIXB7SArA/3aXjsJf0Kk92Mmd0e3hBkvD
L50Zh8rcZpenCmS5/bw9geyr7aQpTuiamwWTV07+9uR1GmA94paVBsuvXqTziwtaGn0v3ZF9m6zu
7JNYPdmm/comve2nIks7N6nPbIvaed2R1w9NDH3FdN/Tl9DcsfnKjGfaGgmIxRP4YS4FtawbP1uR
Y7K1RaqOqoq4IZgV8Csasvv54m8JXx6MW7RAZBckNg/E/k2VOtCWxzMhvKGUvNoTpMC7DtEGR+2h
Uka2r+3L1XapiQIbbWzqQoPJKC3x3eMq4TH7L/8TcUfTRk7nV8lvgpnjf7t0GpkuET1SHvXiO19v
8l0tupMBH4LtWPtPZ2LnUiif0oeZJZ2MVZhHg0FRRXA01T2Twfm8WWg26CSijy9OU6nmXkK6mrqB
dy971QAdTVwPt2XyrVXssatcnFmp0lmyD3WHp8vQQHKoc7Rx96XmPySDC0QPapGodvKZXcXvvn7h
o8J+rplKA82M1/OjEO89z1KhZ7BL9eQYgcqS0F3jMTF6jtBtZe+qyARktaXAiA78FOgE2HZpcFph
bt8PhVIEpXkdFvJwoY4ntUEWvYH8n59c3jQJeJwtU91tyOAHAWSxKn5YwGEs0m4UEIMJVguwW3OC
4MIy/Tx+vXAGwZzeln6NWesoeO9V5v2Svbxs+A2xKvZQdggjEnSDniDVY/r1cQLKGi+dtUOVE3pu
xvxQzcNtm7AaNgCYGEVK3dK5KkNTDN7SE4kLGyyv3js0zLSwNFv0YE4JtPeaMh+23QeEm8owZSkm
cpniJylYcReP7aENUtJ8q+uA4/YYMX+1fxtr4bcskjJiiJjf6zb+iYjGWfPvQtLEG89kwBo/VCOu
/9TckswNk2AqYmaORaS4AI4Z+Q6AHluotna81S+wQn2F2IH50J+wWhKgo/lnqwe/RmIZFq6pc7Zu
Ulg13tT4l2AtNjjzy0xfB3rCGiTyaWhQBFnOtEdwqVFUAgt03x0MoHc5BBdaZQKOFbNj218MgU3g
kiPWeBnxsruhSr1O/ifp1bnbDB3J9DBBiNGr/JqkpdrlW+z+R2COpsIwNz7KqJ5aZs9znooq+rTn
NLtNkYo6Me6Ep07TUxLW0eW8bWxeYNZH8ADqUZYotAI4H5jyaT4kg2fJVqlE86OT67e2K07seJFT
+YYpJfCcf+qJey+D9sbwswZthfSWRgzV5cG15pLDFxn9onTT79brsJW2gDKgMIAzLR0I+A5dQupw
GYQekSM6a3nzamJ/tAvvXiRY/bu/obHZEqUukZeczDYAa5Wtr0B4ucKT2SW6U+t+ca5LaQfsmi+1
VtVKRwfY4HLIE27cP91j/23SnYb3/pkCfgPViEGB9R9x4bBvAudqMamtWzj8AAX3Q8wLyjaBIoYK
VWhZWdxEUXUrsEtL2vwEVQ0F2RyIpOkEVKJMtt1ttbykqvuHN6eArf8LccrcSPu/7caC0rkL0Noc
k5NzvyXhG2EvOyvZM6hg0Fy8a/f/4p0RwLmaiK28Eh5kSmO8t7dXTa0m34JIHijC6yOlg2yYKkPN
ivF3DU7EDm+/wYScWFmUV/BDjTT36CbynT8+4G84ezKdCnaCohAuF7jshERMX03mlDto6vl/JArD
x/cCJs7UMtI+b5OcRyL8aafQaqkfKUF8U3e9h7UQ3jrSNkT/rHqSxiNZt0qqm/4NIvrqxXLe+wCJ
g11V4OCqZCgY0/JjuXur4REa8xrpBg+don5qBygicTUBnC5LEQNUYzD8NGgA7y+donZKMQjwYduZ
cP2hm+twC1VjUHQatiK/ZxxILnlf29mqsnOfbAfOoAFhd832Z9eB7suBb9t8PpLFQcG5yt+GDRJW
B4tlIgR8GRHnOEY7jVFpqFu6XQ2VBFDT5MWJ9oGWbPKB65haoKwalkZz/IPPhC0hgojehXSOx0yW
BAm7gE5OY37A/roYFPD9iy9ZPuGpLDEHQfPzzTiuAB9cBbRK5pRq5GmzV3leaNWEP7tlSMirDfHd
CTSF7X6mpGXb3YoFOAqiQfQwEb9bNHZIBk92p04fCvAxUn+14cUU79Vl+JEXFSZVO6SxAD+8qLT8
rLhFRMpgsQRiihVJ+n6Kk5dtj37sxMZ+m99sLEJLJkQ+0bDA+/ln340tcTEOEl2i56H1DOiZCLSi
QVVxS7Y5TCMMTbrWEnQbxiIV+iPF00cmBjWUelbOkdLOnJX4JTRmAG+WPe+a25cinanCPh+hu786
LuALURRuCKX+Bya7JqHvBhsIaVbwN181mpcqx0OCK+TAy/lVVrOwnYcYmA1mCwjaiGTLb+De0gES
8WrwS31+ZKc44CtTHIC0xCZ0MzjW6ODowkIkP69QyJQev2OB6Lfse9g1Ch2TbeBLO7aUXmXwTUsn
U0xfYo20HeZMDZTG1b5wf0bhnEYRCdn37s+ubxkWUIWrbMuWQdib3kWegGgBXzOkvsZIELPQDW/z
erFdx16JPdx5fr0bhUJeBSq1LQnVKk+JNYYZl3UjJNZ/Kqgsc6ci84wWv9JYAeQbbPWB2jqgqSgE
sHnfvo3qujdfOySwj+z4zOsAswi3kvFgdDTPyWA8VNWxF/nNp1VwFrcbhd+YCZiAW2xtDJutQ51N
XQRv9+7Lex6IyFmm7KHcq3AHOZsQ4QBCyqEzClcTTBO/tiS1nfMJBeMGu6eHfR5v5Ufjdht7m0s8
NoKM3Pv0kUrL0hoMliVk59R1RsuFDC+QSClZnJkFA6/Fb8/oG/9NNaU0pxoJ6EgvBjyO+OEn7HW6
QFrO8but43HkmEzrBx4AgRtsPL84wDBbWqS9j6lQyua3vksx6XRwxE8qGB2KZN3fJ2nKbzY6wVJb
1HWfJ4+m/iaXKc6As6suaN/8bUbk7XmNMxla9yKjAubIcb5pNqnyQ31D/pYPCecursmrAJNy5cQT
P0UHK0UUsZH4OT3cf5n7LtdrTGmlphCM8G95Ct7kdG9fgiKxVTLO0a1sbcdjw2jTi8zb+STy2tA1
Z7ef11nCJ6I3qinxNh3HWs4BLo/9rbgbR+jbKUALpYhd04/8PaTUOpE/71jnEAxJBaTapiqixrp8
5qrGGa9oEQc8i7TT3kc9cj6Qa8hU6iP5nIwBWQGYoLjTlPW9og0oMI9rz7uTEgC5U9qSLnx2ZjJ1
Wx7OEoCmBzbudfDpDfyC3+8XZQ2P5jiapFxiyIrhN94BsGxGc+5lE90o2WNXeqdqzAPV1qbIiGER
BrfgnA+6bkY+iMgaj6V0z803PN7UbH/2DOXMLe0ozUTTcQmd51uzLZN0RptsSJlrkup/SuMTt0Ud
FqpASo0OqA9RCj0OIPYf+TQy2po+ViHtKMY93x/44NB92hzv8AeyuXY2ThQ7Gd4qZ9mldOwnCGB7
r6LBF7yHbJrJDdWpYldZUpjZlJaPDP21KfWkBquS8M59+gR/0fs2C4liHDROv+Cka7dUZx7XVlh8
lg0Nlc5Cn3KXkFxKgia4IpqUxVNIVcFVnT2UE4TcxEXeU6M2P00RKtJ3tSiwk/86ynj3pk5V0POZ
OwvFcKV5acR/tOJFnHDKYYIScGoUblWytURvcl8F09GLB+Gab+1po7ZHpMwMdLuMVVgOYoOiRDeJ
bryoyUmyAvAraMEX12ib6NCzTEJAmkyQZYTCyFNIcpOPaJV0Bvti7VgrPndP2MLOoN+NQiZTl9/C
nodNM2e5Uztk1eFJ9zyYHkGK34/hlOmSn3ddg7dXZDsCdHUY9YSq/JTeMDroco+TgOLeJuDMMOWu
+3jSWvu9TWzHREAXH1LwmgzMCcXZwpSPUd2xjnYoAlRFtjNX0pkSw6IkV5kofzL3oWT9W/ZAo/sC
/fnPPgcnGxfEP6rzv7wokX+YQoA5Yxb3uAZ0uPnYSBZYudCcaDU78h/aBVBRdTaApLwS9hlEmOuM
5kwRTGc7opwLvHCmSY+2T85n95Iefl32ICF6r+VhUj2oGL0DFdJv+JX6prWE/7HolilnkP7Ifm5c
mli7z81ZFKmj/Kr9OK63jO3EIW8/SmHzYO0F/XqBuavuO/Dw15WYgLFK7c5Wu0f75nWYVwbhhWIk
S9SG6F/woLC2e4a/2urKas2TAEslLHa/sa4A3NhIr8BHUfjK0NJfiO9Aj2486Y9++9vzWOvZJpNp
+JPlhSoetNHMXhin7XnU7DP9BUx2ACfP1V4sAFdSWiBsYi0dm9hpPz+IWhakRh6/FDdMEk5GHtJj
zRfYz92L8DyxH2hfpcfV1iYO4a8oYaSeqES0it9vmejS/fBnukKRt+KjgpACYZI7Ooft76NJgs7I
5iI/tEyLeFCy6nfYCspL+OrY/3s+U4U1FBDgNo7oU+LpbR5r24aVvraWxG5QSPzd+IJo3s8SAQgp
IT1NUFRPyRe8b/vqytRM/DnF0KfbZDieyM91FVAyc5w1Up2Xy5+cDS+MAjQDkaW+4Vf+BwgpDkiY
e/h1Qm6AKo7f8A4nIjsOe5ip133jIK+ZisdVeSjL2qu69z9a3wow0TglrbadzIWDf32yBpAMuCNs
gTXHxZ16Zp1GayCO4cRPbP9MwhrlAQFArnMHai59o/DPhI4eCa3wHkyTiEblqrY2tUjx+LAeuF2R
jrAu/FuW8AxlfTIxOXkIJW1Tt6GJ2F8bRAFDwvnhJYLJ50+xVnRoqaxwg8aQvqf690m4W21hqtqj
i760nTV7z6WM9m0JVh/kQLybbOsUSFxVliVD8cJSL6S010XXkmJh/bjMUmbKNOgKX2LvTgxOmtk8
jVw2NQ5uM2ct9gW9kEDZIUhaFYAQcSw34O+T+wnVrFwAI3yuJuGY7nSWyFqgTymkuMOsL9TcZ84u
h6B9I0L9qdDx1hctHgk1ZFGpdXMV3H9PLd0xBOLWaWMO2OXAzrW7naylUfT2fr1zEbMgU+5uwg/g
lbCtfJQDl3fT5GW2FRV0mjt/a8ZxTT6GyG4UPQInFsBEIUYC3mtUQ/8fxD5+KuwmWxbswabffoeg
l87r4woeIUIKnzCiP9hpnQ8YGT4jMObbWNkb4kDDoC9Oe7TIOT87Be4aZPXV0YQu9wi/kA9Uj3N7
eKwB21yWldZG6TjkD+v3Q/HcNkceF3HFnSDtcBH3vpEe9yZoYFTmuqhAOc6Jaq3NxHG4L7SxMTik
vy+hqtBAKg3865YqXk13f0f9EelAsQuBiItxPi3AHvZAmChy4MaaXKfRuDPlebBeRB5qKFtJS3fB
zFW8uEJxJMiYDb3EEkPbVohZu39ubptBhLWn3cDJqa7ytSyRCnwpcI6Y+JcOzCiwMJ6UYbbPyiYn
AI/FW1yxE/WQ4jUg2nfAyC9praFUgYYxmA3tbdxpaiiqMKc6C6OGMXtjcM/D1zyOpFgtj2kzJDdg
0oNlM8hgK4xOHeLwA4Rv3iAe0DKwh2xI2XrHMDQyJkWCAuEZUdqicalPRICZ8LkD9u6XwoehA9vU
L0cSLb+cfYKly4tPzMQ2Hb4T2b+qxMBddCT7WZz80mR88nHazEhoEVMjaPCj7WMpYPoHVU54KYkk
hY4n7Z3dYITJHVkj3eLVm5fvnMLpPLLj3X8kTLqS3u7Kh2OfbC+Bk0gRntbI4xsVi52CGvQt+Qcr
yMuCrBjiAzLPs8W6O0NTSJe+ZjYYgEusgci4ctxNcDSbh7SQGpJJCOu5Nkb76q68gmwIFc+w/m2Y
tb9rEnTVIVO+zPIXMLRWQpAGNuNO7px7uF3gRlreMBtG0Lj3a//cupw8eVtfsKEpbCBMa2Rjy53z
aDiOqoZnKgGCHSNJYXFT9lFKRZpt4s51b9mT6BX5QOGj59cAlzi3lX9K+GJHHCxqVjAhlwuSoNjC
ZuSuCdv+nHvRW0iCep11W93WSZl1OgNxHpcxQLDRGwT4h8KPhZpUqXrDPWC60POQmf3cVBUzBSp8
/sKEJO5W3oQQqu/Nd0667M9nhxw0NAEbjjlxO/NN50yc7tpra5kkl6jTIZmPWw/W5h1VtWYG6h1i
ZhqvuS7PmhaRbETHvwR0Nn3svdXT+afZy4KUZgeKS9RkT/5v6KBgKq0db/9nAeT3CEnv7jaD/tqH
1yF6AYgBhI0TQVjLRgLs47BsU8tQDak6UJ3e4W+6sBt9EWjuyCiErjF7lm7fx0ZRRIWge8WHqINY
CnKHOV0ytys5de5kP9eJjn2O3TsXU6fIaxOJgyAnobdrqOWcnP2sEDkKhNUMoCq0monWp7dW/CCb
VTEHoBle6icFkUldAoaPCu6RiHnkaId4Sr89qEDg+MQTkvWNHceYdqL13ClCbGe5pmGJFlqHHhZr
AVuoDblYv7MZIZhwkkCynpzLJzOLl2fnMtNuCrAuDswEmfKs+8bH6TnpYfm2dNDKmMi2apuknAZo
zMXEF7yTnkQ6taEmj4jmc4al0icJfnL7jiPJYhdgZoj4mynQq0yib4YtHUN8cA/FMFkFO8C0Uley
/Fdj31fCIvHxaLHyhLwnlAmPVZ6mN9/JfmzO+T5AU8mz/+0IcpDpSGo5Ig6sij0fP8UTfP8zqqBQ
36q/7BXK6l41fiHiN9h548TdB+4qPDEejT2fAbvxEAyAJ7bIWQHKuNe12cFuzFGspnoRONaPFEJ7
Jy1nyG9amUiWhbY4MhWn7TqLQr0lQXVTiMEdeUl8bnPBkMVYv1YZkelU1YnsqatkSmregjRPJri+
Fj09B12lCyovNgecIJYahOidabr5l4BZ2/HyLPELaNDj/BBBUCk9JheLXHy7Q0qs+lZVbQJzZydj
Uq1bQlh5lil3f7Ep8ha6Tm5MTatfWIYhJq4y3LYkazG5EFzO2exh5Abx1RtnM0dVTssEg31+Hb6F
86wL1EY5fk6wZ9HZ/97Kn/h6omLt9DgtEx3y9GuuLVR5wvbs0DJ2N7YizHyZuftYsQV8Qvv87lBd
isnmjjnr1v+IzE/inmE0exdFmDdjt/WoqTFg4t4l9fuv4ZnFIYSGy7d77Gg/n+duvGj9cvTBaVC7
2F2i8Et/Wgg3yA+rkkJuXRc3haro4QLAC4sHE9tIeuFnrZ7Ifui7ccxB6bXHpipkVwtjMAFHvG+U
iGyaCRdHsjbLk4x7dHuJV5NzId8k6Y1B6hUbzDxuO6PKNY5VKoZf1ZJkDrXBUPwJgplHx2+rO2jG
w7Vk9C8VqVoFLCiPtPV2TAzV/TtzFjx8DqcsQERXM+1TdjYFDXe1gafEXrcTNAr4j45V8KK7ShBj
FVyiD/kjDCYhCuCl6o3ESQ52fAMrNwtFntmS5sEwtX0JHJdwY5cVrXoHLMeViOW0JEehcMXpOoKU
5AQN29vfT0xtTZ31cW49uJzHgGbpjqA5PSh5f/7P1n7pIVXyNLjXNxJ+ChJi7Ls/AExoUsZfHUri
iGebwO5cGaCk6bZ7TGDjbSi6yTYgcT+3rWxg1Yi4hmaPr/wrfoUGXWOpEWXhD8F+xSbFYK472Iwk
3NAZXgsxFPs+AkaAwnbPY3Vys9AVwAPR8xMGzDqWM5uyReFHgGdDKk7GliD3qvzLwgb+Z0IUAcZi
cjqzhZsF3oA9C/W8/nbukWRyO7TDIpwJTZH/lP/vOad2D0YAKuogo5yLyCXHprDY0Ii6x3XjtCOV
5sBBl6O2lYodNf0TrJaXWXSQDMfU9NSfQ6sQZDnzOc4jx0MgaUhdiy2p3ILgjP41omBE56S/1T2V
jY9BAhIiz8bhCqtd7qX5czDMsClAKijkfPM5Vv+tokaxIps2F2IioBYSptJF1u4tKqgYaD0cb+6N
gxnQglFR7D1ZQuw5JH2FP9I0vW8+3nqjHLJCWlsQSTmSiLem7vbowoEaBuNMSA3O63zQyOYDzJDH
o9lx9djJr0Hpz85nFzVrqdCmlnM+yWveajMkaqEvxO7P3Q8Lr6eXnCGgSlZXV4bs2v13qeNUheMX
aYPWwO2H/BZKZvQZUrRiTUjcSQh6ImQwDti26BqhqdDDEgKHiE08L8oPLMj2qitya6M7xeDHJmP2
hqDabdGXBwRAJ7V+f8sFHG6RdliYNTwqTxYnVv8GR0UdyRgf58C19YPpLr8Zh2XeJCbxbC1HReCW
gu3WuebuKg1kh0jSbZGtYvT+0V8TgUpP00rrrHKphikrOGDYm5GPT/PdWbwa2ZMNPe0z7pNIeQ9Q
PBFSfCdJMSaRvQ0Ilo7/Fagk+5B3DIUq2u8heM4Jp6y78YM1ZI46a3u1IW43pzRwb2ipWifGz3ib
4Pi/iq1INBDigOOi3Xuqjbt04uW2anJFdqQw6WH65SWR183th77/nqTDZFjccfvfdENSJaDFuemb
yVUXbiZIRQ6HNWKsk9+u6si/maEo8vPWG4hfkRz27Yz+Zrdo3re0kN5Dgjf7unHEjtm6YqdcW2hY
RKr/OH9IioNswtwGMKW5TdDK47CR/ueNFKtbYZMr9RugFnEqKNkJ30Tr8UwtJyhyfjnqYiZwB9IZ
t9tiFyKLiBOBYbNlu54rzX0VT6FaHUaUuLl8F5YHkzC25FWCqKPi01YS6ZhM1PQoAuji9PtdO6J0
39F/hwT023FV9+W9OLRHKZEWcF1t9CxMDnbgypVCnEljAMdG3lKXaPS3TxYQbSfcoy2IL07NtWcj
7/0Z8rt07nROALD++W0h+quIU2iH2OpqVqWDoc4T9CaFemR4e8SENG+5V7ba8VKtb3PeG2Xj9BYh
vLG3JMiGcNofeMza9lB8RCmdfi0xnHTuuP+INSfI8feB6sJmuYA4ia2l6YEhYKw9h7WmhbzIs/CF
Y4sBrYjeTFZRKfsk9GOaEQK+BoV5Yv7X+0Ne1UC7mm5UtK4IMkbldyRKJhYPJsNLBfejw/nSqo0Y
RqPQT/iSOgaUIfGR3ddvjCa7z83Oc5zsOvddaZja34jQolGWaJ7rnBOhhgtQvkD13ydzJ8LP+quV
NaddQ8IbwxK6kw6FIWYqb8u2L73yJh0BNZzXmHrSSAyu4HPoqRYc45DZAHYRRiVoMQg9SaDJuUIO
di4XqZFGWPMNmU2Ra2g8J08WNMAYqyIz1uletkB//FG1EHzpuANbZ06OJWVogRS51MvHCGbZrr4P
bHaA8+4mepLGNwwnGGy/MTnwHh+b/cluINctaJkLmK5seVQcpSZBKdecF+L0F38oHCjjGG/PMV/G
gSFwfT1ltMO6+TbFLYz4B/DijZXbH/7aLhyUAJZgKXWo5G5vr0EmkLKqggc8wuePoCRVdUGOmZJu
6V7o5O0IzPJlvivU67gFlx0LPDIOE6odOPJ07Gs2a1ZIhchoXcHpOi85s7kdJQwuw9JdpdfDGEWL
SebH7Rwi6IMTu3dLGvVz5/TytgiTs8q11vEwrl7BmxKSW4x+mw+wBHnfOFbxFLpuezd3IJf9x/nx
wmUfWkRLC+HVprn7uls4/ruZtq4PD6K5pCLZ3SDGhYNK6xS8NIcz3+z6CAtyKk3u9bibvma23P1B
I3WDBn56Km9M3xvKHPN+6o+fk/IBEwynbSlX+xt6k++KrsSw5g3qvNg1eAhs1FyisLJqGdPaLJoI
irwVgWEqVVKPinldlsH8fjsD6FS/a6XamkR0SsRTqLVX0CJ5KDj7vNWgoq7nYvGuj9wyUOi3sa4W
LJEDxAKjjH369zlUvI13Yal2PZGPETQGUYaP5JyUrhsPJ5GDK+6b9kmCZw3lnVMQX+jhWtkZIcbK
3cN1//HTHQ9jeWDAopLsK99MyxyGlUu0l9S3EY5g/ZuOBTlbcBGhaM4AVBuYUBilqWgwBOUsX/ug
zYtV0UNB/pKIVZJzKNMcjq5FMDDRRlzy00ZdjMn2oVP5k5CcE0mceO2ZNNbaIeYqYlm52fKldwd2
5MbXQPTnAgPngnFqRq5maxjCZCqmTlT3K2Q2JEvgd/apBqvvq69RupM/LcqxjHxbsztbQWypK2vd
ivbbazDit585CrzLQg8UQytpRxUOyy5wjFmgZlNiAz+ecz1J5hO+Y7S6RK2csmc3yPb+xbM/B3EE
rnmXmhQQEjWBf4cJA7aAzrfjA8sBO8sySXP/4SIGG7STWcZqq/FC1UPsJ6EOJuBC1xM6lWj0mv3r
+TpG8zAQPsZ5ezTedpVfYWV30U+wDwI0OjnDLmdwE21bHanNFs9tPTLYzk6YrGC6Hu2sw2yg8leh
3tN1M8lwE+hhUrexqlNM2CnMU/NgsCOqK9K/lxs+r74w/2/QJlbqKBrBKwU/PfbIH/O0Xk6NfCZP
ez7vUe1uzBSAaJvPwFIFvxsT8eODUJUCUxXBGyO6J9xQCPEQ2mX1dPIxciZwa/lUJIEzUK6daGFV
fRyuRJHnyLiTer61MFygvbqYqMu31XlnxjvosN2EUPvxen5iOe3/+fUlxZ8TmTgJW8T5Ym6VgMVs
sTxgSigYOzKqYHOiBfxd6gy0PBWXVuMvHRhpeuilSFD/ZycoHkVHb7v+E0ED1G13lH6MxoGaV4AN
75HU72UlXmYLtp6qzEN5G09bQ+onEAi7yEvXVrKB4P4DVRgZGJuzZTfa0oPaoL9DNNWsXidwo6kQ
ypIpFykRyj0Ii0EvFN/LlWd3tU5jrOYCilriMEhPF92b8xBM5lEIEiKcJSKCZQrU9UtdrmGY11u/
rfZ+hTE+pDSaNXDnGpHuAF+BQ/GoAIq3vS2ZT1Q/Mvnpt7FDcIIJXwJAvQc0j9Lv+/C71nf6EL/O
1xDAt0dM5C+SKrNu/5Zjx1aI9hBjd0AzksI892V0FzDD8C/LOJJ8z02cvV3XxLUlAt6RuKDXK+sK
kiQD456m1VkE2PaP6BzzOtAvxLXf8L24xFynKXpAE/EZ3171NeU0PjWRf9vZ5RaSU2jKFUBtP9na
kit0Hc0IZVmWIzh9ABH2uMEcGBChOarw7scvp5co/dYsq94Yp1nOJQzQI4LgsYpaoy5GFQsaMNg2
A8EGlRyZd75NA7WpkDv+U2XDuBsDHZ9AzBrJ0nCuSOKNb5qPkwyPHHd0rLQh0jk99agquAgCqzin
+8EeQWXrFrEXM0evLtKoTqQU02ID4WLn1U+5yVZXCvuqU2nvd3ebbsKpOtyG+tz3YQavzw8XHquU
My4aJSiwkfnzcJZY8Y1q9napy479BgN2DSmrUWM4B697FeRSmtPMTw+sJm9vUJSUTkleo2cgzijr
5nvYDysmwqq8ao2315OHZz4Auho9zQJGrZORQMRni7uOX3NSeeefUtGsYw+EuO6U4pKX5cM8LvP/
SJvzZMzXSHOt0btkn/D6cS34uRzPfPMirOanDLqBcUcrq16EjIDuVSeLr6Qhw4XS0K9tcCG4swpt
Nc+JEREUhlRaCFHbREOVKeDbkCWRrS62hsbvXS9Pinj5tEZve9Hp/29lKR/EN7b6Wn52d9g/WaHX
EOjMSHgy4B8ibbDG+mLJQSf4LM7klsii8CymtKm+NZ+GOSWKGUzDwWyXPeEG14UaIWfyVZRtnmU/
vMkU8mqwuOHAPmutUJm5pCC2JQURGcUmg3AP3LfpygFYQlwoxVdAwUXh53Qv7ECZwhKQJFVSGeC7
9/ICKlC/K65apTSDXJAdDB7Rb5VBiGn4VabgBz4QcbmptFNr7i8SMQ9CHanmcLvof/jHLqxf3AXl
eXUCpmLD0/R9tko4ghfumXZfyAd6EjSg1qceIQkdtxIsFtFz1C/dcsSU0eiv9MG5lf4cc8KwmniV
8EDheo+9j68LDXcJF5Cb9MsJZaUFbUVvoj4OnTn2OabGFCFQHnTxSToiWrIG5omIlIpKzgacHTjz
c8hoGGXqNEN2tWz/iC86p5fIDFrmtbz4uvntxg5v0r8awvXlnKHwkwscAiWdjQxbto1pil4W8Ff6
XAUZeQ6sdh/4BRT39zGcxadF2SQRNpkx1Fy12zbF+e4qPRiNJZM6VqW/U7MSvplbEPzUrPJGQ8ef
CIb12W6PqsGbnXtXFAtCVyE6fSFZlHgrw/Fmo0N1ReihsS945n0o6EOg+tzri5jdQRvELwkkmacB
XF5g6DSbjQz4jMGeHe/OTZkpLu1cD9mLqCaRfUlhtZJxAgIruKbuU8l/A1ZxbHZtOV8AEzoF96fG
ashtl8hak4gyap0bQcryQFrcRXBAyD+UlactkFtbj1SVqqnGhZUl3GlH5e7BwFMd96WWtr9Ar/HU
FrmIDnfi153a0foOrfZe8ECLUJn1IgK/hXuzkjqM9Znmd+6NOryX5W2gycF4XLJ7KMJTeUcGih4T
V1lOwCzGpaLTYi1ZXv4rS2zBpv9FIY1j1+kmKGAMoOQ0qNtTpeiG4mnQ3kc8XG0/jah4rYRZj84N
Mm6GKJBZDH4xrzKEAW3RvO14BjG4eqNPcD4hA6tV8HPv9eApObPI0bTDlN6XK/RMUNrYejePQYBV
XiEuXmerSITwvDNXbGcnyt19su3iF00OFM2fem5RRBmyp4otGxTC+CDxyt4PsxakEPdXAr/eDl1j
fh0iqhWyDblphADy98icdKVC1roTb6EAImXk5N9DGJ/NmGOshF2ifHXjg17fZmZOLgjzDc5zb5s8
Zyr+rh8ZAQ3p0TpLbmZhI7naMgUkqtiruyrpwE9FWy+EGCU0AeLgjU7+r7d7h6TWhb+bWPLw88mn
xO1Jo//fGy+ni3ULfjeqHR+qR5L7cDSbGPW+U94lAGPAPkk6mkF2+zOVs+oUvceS/9WAhhISs7iF
e6jJEEhuoN9tFAnspcZroryZsAfKOObT5qCPqpGKNKHZPcwtDN/HcPJVnEl1yyw4sH//UAHzPcdI
sws6zhMINs6UPTs/JPDwVVdodaVxMDG0qpLMsuZY5SLt5aE/oNHLzmx/H1HekGjOUWBXzCta3E8x
0E3A/iSsMpjyK5V9D+NfKL5mYP0I5TTgIjm/o3e9J9lfAE7iwhBS4AcSKDDP7cUCxbl61qmowOKN
ZGrlcJ/uDciYgef+LtJxyfcbNZleyhqShRYQnxe7DBqoSzuqk3aPhTuBoOUEAXqGBAwFKhk1Wdew
QLuq+gxapv9gcK9AZhAZwiRLnnd0JYcpnpRYWP1cUnzo5Oh7X5O9I/khPeEFZy2AFjTVio79/A0g
HxGzULpukd3C4HPCCqkYsPnusGduiBWwjtTMvTk2UZtQHqXfJtvlCDjSsWTm7VzM6PjG7XX1/5mj
AEp+1D48UCPhGA9hNd3L6UHcGPZDmt7WKzA/dDa5lWl3xv4qbg89zOyyzenTKgLH32L3wD5L3vOf
DorL86BjyLrrJHoZnLOCyY9Wx2Se4scK0H/CCLS4sPLnO9w5SK6lYuddCdDjmNz8tPHJ486QHpp8
+dknkaBLxw89A9ADz7dkUqz7by8S1OFjJ1MXMs5L4/QqLOi8EYMJIWpDq5jYPec1Hs0wzp1P2tT0
jvqZw8uQvx/8HMFm5e5TghxdteC6OJRVQeJwnM+z5ndAMxrXo7Hjyfm3m3c+q1QjGw+8XGVBKC0K
9uFkvhsrA/kLWrVhVYm8/QV0EKp/cNFkurdfiEEy1+wFcrMWwEMKl5VWA0oN9MMTQda6tPsWmH1L
TshtTeAG1oaJbahqq1fXRcQyHajevgoNnoJVjErZNJn0DJwtoTBXXj23lppXkH/LmDtm94jw+FiP
6Pal6lL4NrFoPJIsQejAazTODTaUmn/hHp/ZV6eZTU+Bs95cLaxxa27iKkcLvHCLVBtYZSqoF9gC
GMpuJGwPptan/yeo5t9wC9zD20j01r+fjN3vvYBk3K23pdGGJUcfBFI6oYVgjuqNIdLYLS9j/Mqc
N+MTuUIhH7VHhG3lygTKzhMNPmRnnYu8RrWfWGQTMdxUHLOVKPsR950NAFU4HAEUAFK0X+3TsmJZ
NrscbUsCR5aSK/mFgwPaPxCJX+CkiZCllNbM2bAxJwJBJpQ2qG5mctwJUmybY/r0rPg+WXSB2vfn
3E6/5fNN6TI1RhY5jlN8Ql/54BXmGr4tRaEMKSztiT5mqM7aVxApw9hRS6307RVzoK4Pvh/qNKnR
2Q5PdmWBbm6ZFhhpLhGxn7y6KcuedgNfujMvuahUQEEvcTw1jdV5PdrjdOQDaBV/YinjFXijIIog
+UdmTYOMUSidS4ApdoI28QeIXkEV+2z5Xat1lGfZT4y/C8YzJtaKKi/QRBmc40r+opwJbR6MFrQ2
yfQDh8AyNx5extvEEUtnHbHyPzqo8R3UmCXwJrpDsq4gLf6YxO3MXB8ug6/IN0thbc4khf72m6Ca
qbXzJ/Vcv4VyCR84spyFGSR2Y61KoLU58weNkWvsKXr7RJTm5wuaJsrwhQcwEkUa5dtOFgf94c0B
+nwcqWAdYnIsXHovO0jQgrVE+wRp3vId78yjtPs7B7cOW99PeVu16MT0Fy68VgxMZ9I51AoP51Ul
U+BsdulDEhppkPay8PlfOyt7EgwxkSNFiYG3fMvJQv/98llf3FGDqq7lkArPI2jT4WY/F5nZUpM2
klZCqv5gWXX8Kbhb3Lu8ybtoMGfRZbkNoI+341EYE/apiucft/ZfFi/cQQfro8ltL1/2pbjIFIwA
3ThJjm34fnzbrlEGUP3MEvHif1amwnuCUstG2FmC09TcTTdIl6FDwjjD625TbqlIqAl3QJrRGbPv
ylPHvdJI9XQcr3rWrg1/CiLJ9+cES57FgwyC4BYUfYupv8Ix+s1K5AOlWlXYEjAn8gQ+NKTJG2Z6
gwHNNq+fuI5L+QOxhFTu/oxF4K9tbjFSQWwDQ42H0RIrNTIyLMmK/d/wyKrNS8zKJe2gzZQAPiFr
y62WmMvMtB1Qr32hIClOlVYK65MYczIMKzo+1wNfyoVqHE0revJMKOr83lYYzqNk2TqvCHVwl4PA
lwirmKM80tEoYzbhebM0O81MK6xHzJ2R8Pyn3C8EzHu71iHaHEObz7Q3S6g8hn2WXEAPi6YT4K8x
ycUEaCCu2lbBHTPEfx6Pw2vyn/IqTn0m33OVig0Z+ODowNzHertp2FwG4JHb8taSEA5amS1yZPnG
NoBGQf8TloPUGTful3PVxLTc2FNyvki6JtZa84U1dJh5pBUHQ1YCHO+fnA4BdM88IlMztMqaLu09
qjfXnlCN2IWYFR38L+NiUZaykIDuG7CFd3i7uI0Hq+fnaiB4J0gI896cj+QKh2Rmj/+6cFK8lodr
8T8Q4p1ya46r8FOILqf06eUqpJ7GNSWm+K6ZXz/PwosDjNk5kyD59suNS4kaYOHUd5g2EQXiV5QU
JR/YUcBNc+LHQBz57OcE1NtKk/MGdWSaruXimDyrC0VUX5a6/q4XUVApSrt+JitLfJKS7hBwvP8S
v1aTRcx/U+qJpQyD/jmnKfLwrLNFQJLLIYBKH4yRPeZU29AtK+3mnf1/nkkozcSD/67jGjg/S67u
o9HSt9NemTIvEHQDqRky0ktomn38nrrbDDkvNx/8eraj1aBQpYaO3QBPc6M6Y3NzD9T2bhJVZduS
JMQwI8RVadYI6gmayfi4+2Hx6Q7KHS/lBSY/cmd/pr29fw7hlDp0UG4Kdap88VuNDemOrVXb1OQm
wIOi0TnrWg32jH9WN1wIZIQyq0DJWLQ4CeJDrRPkhd/gxPADfyXg4xP0uGOAFfA+LNZIfvg7c4GE
ql3YVpFbr5c8QPN5aAYOA4zI2Cqu5PGI1uKLqdkVgyxRxlEkk4YeFMx+jqrAVUTkOiOF4Hj52kbI
KbBClHVJSZVUXbGRtCcjAdwhtHZ4Mt9du2heGE3wiI2LAUhSn2RINo6f4tngq3IteJNPQBL026se
zktBBFcsuXiDzzHl2Eri24DOxiz/1djLraKPkIfKAjxcZ4p4bcnXhm7YjMILCUQbZ2o1uKA6uPi3
Copve74ycOy6Yi4++0X1yxeTkdDyd9lXhrfc3+XbkKuDU0WmaxUjrVHFNlwLjMazEYVzzpghpNS4
9NaFOPndB734u+IsDBE+xqHyCw7p6N4k4tIalAMCpUrLEp6dBYN3It+xIf15hsVZTSbR22E7hrc3
r3H5DsK2OWhbhnwxDJ1QCpUVZ7IeuHpYdAv0X9xCMz0qsYv/d3EaCZ4bV+3tEvgCJjpyvnjSzyqX
aNHusiGxCdTYba3nLV+UcUG0Z1yfR+egaoikIYLTO/28QDHy5vvzSxvXuoDV4kgvRdoezb9kdM/D
ajwnbjHSmZYHadvx/55dqnRxZTyZo/yfGxMRcL6+EY48A6gkEW9JbSPSUpSmsZ0vmHdybE2VP6b6
2FPs1EjzzvTqgn5OiEMzDYEMKxkDhV+eHLw22pcWPT3qwMb1mRZJHQCDup19VKcUj/vb4ZRjzse/
vxkQOLaiYq1+ki3RJI/RR8FIwjfJk/cj832ZoORW1nNy5oS1YzwAVzDZnUOCv14sH6qXX95W843z
VYqIcGd5kl2QTEJjK42+75HGZbBtN+UisaKLepEubHr4Pu19tUSj1E32szxtYQb6Zlv1lPWso98Q
V3rVFTGT40HQ9IgWKC9P/OjxA7bwVzueHNpVbUCrArOSZLd/NQZp3AxSsx6I2yvDbPRF7bABu2M1
7E6eIDp/KEglptQKturJt55YuRltLu9ZWY1mXMZhksNarwgsWTf4Av55d/iiQNXPmfW9T5kriKxp
swry1epGnNDUF0SXoMBnhvgTdjGnevhAcqwKLzyf/T5ngEdYeFuo4J/AWzTg/eZPaj90Oe/SozS2
O3vn9MFeB7FvXMmpDx9ilq/QFX0pgBYsGatdX2wFuLuX0eWnYeivK9oHqGRbQrEpNseHFSdjIKjT
QLJSTt2xgHU4WMzlp4QWF0UKc3/fU7O6x3zxvvQw0eGiJJ8iovaupWjy3jlviE95yCS+FZAso+au
5Khh1SouiKmJutUGhT6EA9YPJwH+iNx6J2bMIxhKhlItaWJCyIubJ4elYIQQLH65zHGxemFNAWAx
s/jhoWMqggkAX5Q/xNseaFm4sUQ4JknIYIMsQ+5S+/WcimL2OjFU0xqhI0w/9xu81pWtQGs6FuM5
rLY4q6ilmVFndgBJ1a6fGvgSxvPgWnGLSatMbOL82CixHzKqaYI1i63i4MWflZ+feHuh/e+zpoFk
GDUrEpOd3hoQI7ykpVrh6mzK3+Ip/8XY1JjSZbPwfVGF0tvRP4/U0EBetk1UmlgaafDdz1i0SFrV
pWfAOniEDLIHUxd4kmQ7ZiI7losk7R7DP8vgx05fp0FXUjLNcmZbmTRpB1sCgq5ChRflhEw5e6tz
LQzJw2RoUrVMSMLGwfTft2T/SRHCXjlX9bhjL1AOYi57PHXmn7YYqjLeYorMKmOezWeLt4HyTkcQ
G8nK5gbd6HwmbmRNFvJ3ZiLMSPyMdyivUwjsL3jJyfpO9w3JOGsM0w2KZWATkhqueLtfPHUwRYPE
iNApTnj/Ul1T91g8VI/XEdxsG2Y3ZbK8m0BxmQDbHA06PSuLmhqfMu1h01XiTuHlwVpTiOubq1Eu
T7pd+GtsIaK0AcrPOW+9xxbb4M7y5OZobbAqHuz2zG2iBdsDq+H8QjvPoW7sU1E9tuiqLkLOL409
f8tybdZiI4bjaW9D3Eg1FwnA21VhXJLALDwEeS/TRP7wOUcFTElh0cQnK86tuAy7xohcKgOTF/9s
Bh6aQu+QkuxZo1ppWL14MSPdCMERYjKUgkAZtAh5tI0LP6I0CRYHhfupYz0tE9s4CrUHx6PTkuu6
knftiJ7kNSQX9Uw3/dbNfdm0lK1EjubvjDm1YTpwqk60I7RNKBnlGg3Xpsxcsm+lvDSsNpHszUbP
dMJwTFvIjXhSriDXKldc9swVLq50SKpiIyDj/DpeA2aEUZmXKeaaj0SqK6W1Ij/gw19KfnTOrGn5
s9Vo76KzZC3vMm8DCm/RDUBYv360wj8m1FGn286lAthbYWpjCpDdHoFntTF8+dAlprd1p/+E+j3o
iVIb08I4hRT8M4yxHy5zXSCUiM7eblLbziIlZMMjLrGxP+ccJOU7H/mjbS+ulrveFKX9V1JeK9Bx
e95wzWPsVop6xe+LpbSSipiNZ8wfSAwgGrguJHB0WX86j+Rd3DBmWFBFZgLPHxF50wXpkbyHbe4g
3Dkq+3T9xI79U3J0kEPvhZaeri9fobFkETz6KjxM2svY1PJaCGTHPw/f63Tt18QuGvoRfyo7zZMb
XS4OL3HVRzln8ERyxKjsSLiv9Ig848TYw6NqFPqmqkrBd5VrncjIWPa+F9NOz1kpfhU8bnzqLdo5
L6hZUQtpqXLUfVbQXJDOa62/2G8aNYg7i27c9b+3P1eAU8Gju5f7YaLu/yPiT6bP3d8XxxdRm75P
qpr3kRbif+bKEmCHyW7H94HuQ4LD38bJ9BpWs95JEPGLuXX/zlCUzxzaiXKD3hDPrgWvMgiAC/hz
2IIfOZMq0k/5etr3Dc2U5Ubb7dsw4U92WD38196htdhUYt5GzUgYa/pZj9hKsDh/RNpQ8xmYCKW9
L4aRbs58GBAQSI/q+olR/PilcgEVy/qHddoKhtk3mkhseV0AGlk8dlD62qA1aW1sW/i5voZLAVOn
atswaDR75Y9b0poCIUAUwsQSv6mpyKdg6lyoPZpj9+gYWQn6+Rj/9MGTnd9mQbY46mwO78xFrI2d
huPwteSJVcpXfSFLQa1SuZUGvOaLmqHysa3HaCiiPff51WV3ZreUAc1ITjHBhJ5lfTvud3jb1f08
muqfuZPJlxqAt7sBToxmZ55VULOZ1H1wuDCx4a0HyMDiZTHLaFus3DQ3Fb90bzIhtMIfLYnPbgZI
hciIawkj4sm3NWXfRI017YZNuaVLlCN/WGtzGv9vBhzXBE/rhD4HnJIeuiPLJ0v8WPnjRyvHFKuo
EW0+Uki37VBzEmIxYuhMimviC6j1/ux1pBuQJY2J/u2zVs1XhEztZgCZypJPV/rDH2AW6xvOM3HY
0I5Wn8xPn/KTYdxuY/fRHbX95HoRyZO94tr9JCCmTw47nGxBxa8TSy+IpNDtwefZuE33L5SlEQ/Y
PuSiqwPnQw5N74lwhuN8/jhiI3anbsjyUCtQw9+bRU/EGgKeym5LEgAfm3LKi/+X607/iliVC5eH
jPQqR15FzSXtad2YifKvovR59O0KXTxMe6D/NQ6LNeu2AYDY6SwcogsiCtLMnPQe44GxdtAO9G4f
ZEULgOYEqQtbLJUBKTvXHXjzexUYl/nGaoFDebiOrBnKG3hAxbk/1WqM4PnPgrLc2N6pSl8xI2MI
0ISB4l8L4gcERW50xdEaVh0i4nG3cv1N/F3+67qojYL+qFQOWUVEDRbvr8TSnqx1PKJLOdvgRIsB
zX/RSUPBbwoSVu2vtja9vjg8ipn3+xB1PuwP+ieFXy50h1nYWrY8Ol0bimlkU9jcyQbpwtB8E55X
LR85ivLee8cZ/g9N2s1PFwYwwhm/LT9yEI6C2mBpv5jiAojRYoIXm3sasyiWWL4CZ/PxKa447wTj
Ueoz4GegBxfqRbli6npyjKz6HydltSD5xAqzCL2x7rY+DdHOE3L8CQneQk+mGAZfcLxpoQM5OvPK
j+8KdNAS34u8XbzlVAVNpkncglnwJRDFb2uzi0v6zoa27QSp4zmjUGdSgHkYUROY+cvV9bWcffhA
eLv4MPTOf5Pffn5YkMA5DkMHAUP2FAlRNr32TnkN7YmmhKebhKML0c0CZ2xUIEsfp5Dm9MctupcJ
1e2nCj+XktJKJGxOstsbzSmNycNuIx0Ynbp2vP1zvjtq3w8drln252HCFIItuIFTL6oML7OWmdH9
MbosdLz2BTdxL0uWVHUhhFORUmPnWGTAZ/ElzGrSVVr7cDCcqUBdPIJgjEBFTVxrRb+0ZXhNSuBm
wACp731X0BUdA30cYTlqmJ5CSD5zm3n1WtcTM9ZpPKG3VHH5UCdHB1k4wdvlCNR4KD8aX5rsDQev
z8PTHujXKKCmrw2K8FVOjpyFXrq4kcVluUbaa2ztwxo94BJ5dk7Ex9zZ5HH7Gsyec972MiUPeEQ0
qcGJZ6d0ObZkkVFMZ5hVC3TaWza1HGLk1zhjmiMsBNZMRISUKQDeVdye38aBpMILjJtglSEmhNP3
7gSRCmOh3OWRM1SPCyGmal2BsVRok9SkeicUu0GaMmWNt9M3uQ7WCy+6Imj89xt/e9c+5sGkhkNO
DQCaHFIkQptEOBO9Ny/VBxwgdASj9eGOZcTq9vT0If5HwEXh2c76I/Y1GLKw2bm8uPCYplCXKtMc
PchmfOY7ySspvewzR4AyUrjpIOp1ExCpNw+hbKBSTDLPh/FrX/wRxxzEkcYuAMZGpNnP0UMjHYr2
mL2flDLPLt72WdF6YmZEC15oxNqsL6uHk5YdxBxAIpsRK0Gl4GcKGUY4vMf43zLYL6huhzE9zsjJ
Q3J19mgsgeWV8w4ACSdKjqcxYR0HkJSQbBYkFnFUGIHSaZW1JpLnX8mm2LScrJi8Po3f4fnUnD3S
+91Dhr/YhTuAEgrhAPKi+ZUe5A6VXBvyQWiUELvcJ8lH8G2nVZZSvJXXBTwrZk5CCpw6IcSWCPIY
KbkSwXFWBTDwk9C3gB8+KeqXgjdm+/7TbpOogXkO+S2bh7WONHoudgEQ2ARX8PY0eVvJfeY1iKLr
9nG+0dKFGZQBemLxyqXpEYrWOh2hnPOdsn7hk2Gb5Chz828KheVsRmKzy2M2Aa2Pe/jJBwA+voDA
XiSzNJCvhvKU7eGNMfuM/DYn0FCxZtNmb+YD0UiSFedrsS5wf80gH1udnbj+a4JowdB+XjHBJPfQ
N3xf+7SifjWCCY2r5Nb6nVPTRCRdFnYLYM8CuGsGsiOLIGoI/A5HsNYlTSZj2W7vbJVOcsB3zfA7
cF0Da5nQVq3+eBOu/za/+bRHYq8cvrLzXwSEIkpy/jnVufakQ8Q4QtTlnHhvNV1J8mCWBglfCces
eGmZojq9qvVXykdrRP/JGYkgqrxswxGeME8DpFIS2s+ZtgVBAaqEP/Q5z7AIDQrn34HFTaknlAgp
HYmwYoFs+QZ0Q/iC4yVys9WJvdLZJXLwNa1qH9ysBaHTzZ7swF0Y0rIqYwn0zB4nVz6X+VQp8bPC
WVdQIh+vshOXmaHOVog3QY1nD5LN4aqGIHKI5mA5RS01q4UpPKS1sbwkp2hSbQ03pJfT7ehxSaYm
AT+6Taa+Lx5XaoXtqQPATcqIuvrnByc01tcQBfjNIT/IbPh1S0SpCpYq8B/fqKRsAvdSkEBBtLVA
Bp5FRUExc/fPtKXbY4YcNL//SJuqVKgP0vNm4b+Adj8+2j09cHMGI83rclbnV1iopgfW69en2BeM
bwn9MlSlZiHBomQm2Jx8iVBrT87X5Sgqfl15gnKkC9yI8czASe4FP3hk4ckWEJDIi9tQH/yKiUV4
gtzYVFjim4vYeQl7bkDOfE67p6H7uqBDtpu+lQPlZsR8b7G5jBaeQW12WZACVhOZgqNnf4cz7l05
06Xq9Xco11RnqIkb7AERNwdxXij3gm4lDGb6iCjbkuZknC010E+AWcdhDXe5L5x5NdZ/CD8htslu
rnywhaWYlXDh25mZMKsVUxkQ22u9RGd0EwAKDPRXT2le23Gkzuv1rJOlW7fdT9GbxM9F6IpWFFjP
aPVdtru5fMNUz6o1pha/bz4Y4fburpHfcZnlAmYmLY/bAPsb7JSq5yxiTF+rS8ccoPOA/3O856iG
Ons54IfkQoeR5jMHDUaX2u65DxlLetowqsMG1qy44gDZP1OCY8CfnJohMWIKUQNon1d2wsY7ynQ0
iwW8s445s3n8r7YTg/TczGUVMB3tD8jB/ZEcNqewRL4j7Sklach598wUIQyaNxQcPpQrN1kKVJ+I
7kDRf/kP0Fto05ehyALkO0F0TfCapsZs2gESNuD42VIDOPu0KDvmA3yxtkdfZTissjU/0iq62+nX
1X5RWozDp2CIJ9MO+VgnIkiO+ZTANfm1VXO5wY5DRp2eke5AO78cF86yYQ7nLMnQJKxVzwJMVXlK
F1U4R7fR2My93xyDgz0Ff58DJ1LxkHlWE9gxegbNnLDb9zvPhNkoN5aDAaKYxiluf1xRps7wch4v
KZ4WPFtszN1xofNrEKenotmGAylViVeSCv62qFguijC3ir/xchzUv/dc2+DlnpbzkPAbHW8bx+u4
o+OImBAJut5pIx5lRYYjnZ+ZdNVfT3woe4nMSoKJN5OTobTY/LX8KUMTXSNMntE8Uc6shipkyMwB
UP40/SIfKDHBu4W5RLhkvwuGVjIMNjw2X8fwxgYb2r7VKXqqbWtAE30ctkaaBrF01e7D5+wlPZJy
5ui124LW74YfR/y+RowITE8yZhGPZWSbc5pTLAf34w+/ErgaXI1bVMqYNhom4M3vH6VluSuSnZMA
N9wcOg0xf059txcS76n6rnx0S/+vAXalO4V2mfQJE1zzYXlWjchSMjk3VbB6vJck0kTpnPLR+ZbL
MYpAUMmHtW7D9JLfbC7Aya2ki7ciFlRE6SdSnEqIjFzcScafpivXB54uxplEFbulViKnIK+YqWGW
P583izK4dXDzipq9cEAJrf4OricEQYElpYmPcRy7kEhPDKRTpkPn7iJYXMD1cYEsHkzoiFd3e6WC
PYJvMUWgqQPvrRArNcz86LHNnAWWOYcdOMP8SCj2/NyqvH3MgBNaU9Nhqzhih0Bg1AACVk1pDb1W
KQJrF5TxDIGC7H/51B1CNRblRwExkdd0sS5Y95nd6kBHjz5GT+7wIyvPILQIp1PW64ZIP2g6At1G
5QedN2ITiz4D9VVvD9RFtidrrSmUWgb5gtspONvIaYLj7E8TRVE8xlP92aScsvkVfTkQ/TyaNOqD
RxqyUCMDZwwNK4AdxUgCuq0rVaUua9nRSyejXKiJKDLGxwBTaZbPUvVvx9uWL+wI+Kq9pvCcJNa4
9YLFhj8vuP5AqTIMUsDkplT8dIkzIZftSuwbqCyCMuA7seAcCobrRpECLZbTtzYt+x7Ja4pstYM4
7pPBZspnBbOzSfZjGjTEl2vYC/R8sdIt7KTOKUnZeSSdTRKqUCt+S8DPyYUbgWkp9UNjuiHDjED4
mDU11SiKwE0noWSEKEeUZt6n2gxjbQFBVxuNvn5XZCJQeAd97KLDFpFBoJtUOLF7A8ut2H04UwSV
mw0ImzFlJHwv2DfzPGJwAk9FVsUuG///CzekNevsuGHf8/Z0Tu6bMatmC+XBAQaIt3FAf6pUr0O8
bgED9b1vzKZ2/mzr7ns0VipYahFvhVLy7tgqLMLHnG0jxhzHS1HJEXhQ1cuuKaDSCOxaAFFIdGoO
Nup8bt/5/wZsKJUA34soXbUBH4SuZYu8t790nt/CHIyKGJbZoIQO7apF5Zg/q37HvdzysNDp94RD
8ZguZPmIl4q3IlX/cwxNiKQBIeEgSXRxnXBCi33RVmWNXP3HJJwUz/Da0mpTSbP9oNcB80x6+8uZ
RsQzL6D+biLPosDeJBqjmyBAyHTY4bxeMQD7EDxzBJrN+AM1k2CcRnZRcYwde6LL/U7resTNJezh
UIdxvIz1w4hb3lWfnm+Eyszsu/gcpFL4G7BkS6FoJBY40fM8f1kBSxkvRL+xnwH8a0Ozaye+lgQn
qkjYX63vmDICE+iTXjbNLvNUVQWkx8cN+t8Zv+weRwGzdleAFXTmpfTQchKS17iTdgD6ZwZIo1mc
G72SpogNk3gFIMMg/3BHwQ3EP3fj9T+qq6WYQA5CUml9BoYsgFUVpdeeRju+8lTAuMnoLmyx//UX
1pUbfVSMHbmyBhRkhlrRbZ2r6j/QiPzLwFaj2CiPdmFgEy72vkGBDr/X1m8J1XV6lfYP716iaXwH
ouLtjzKrKNu+aYA74rhfTV/Ew88zbLcX8jIh9wlrrodq0dHQ+0usixbQmJfCDviQAt8txGRUb861
G+5ur2ie2BIMVLomZYQrnY0ACh+Qgr+dglJrMkIQgQQ8A7xTprBOHY4+Y/mZQXX19xw+wOV34V4D
xLJkUv3WQyJz3b8dOrd+Kn8fL10hPByvIUgg+7GKjSTV7K3+u6kMRBOUzmdUqp+Wg8m1zMqJjfD/
/YTpJO61r5C/TG90Q+82NCSW1Zu849obCsyGZBb1icOYN1rUR7obEZBP18lkiIu5GXM2xJc7EGWk
op4P5YZ1K5HJ4XpvRjwLYmhCpkBWjIklj7UqrDXqexd67eT9OGHmGctWWx21r8LsRZeXYsz2EjIM
lijrHcvawEJtCkRXUU4CkCG7G6tY6g42C7p89IzI5W74pFXh+fpY3uBQshHS6HL/pL20Q9+v+n13
n7BrsPvEw0E3xaVtwHIvRUen3MeN9SuGuxsVNAR0K2bKU6q194R19pjRPUcdc4rNevy89Bq26oQt
rM27PkVT3fmIkwSzFRFznpxIOpjg3Y7VHHKefSTUed2BaaG1k0Lp4k0HfCAUCdPdCkgeWsJ3KnDC
ka3ypz1Gx52U2TwI+ua0v/duIe7uJv/YulLcSL5g19bG9qc25wjn+XuwbY+OnctFmiQc2Dtbd5Qa
BM+3rjmPZYUdDwvf/F+WDVyUulY6HQi3yNJ7T316iVQhwT1Zm16rulMSl7XR0P41fc4f0JgEiUVH
KAQ2GgrZsJEPp1MzSwQ9zyvvqbCPXTCQo428plHLkRxal0fVDD8xrJxgqJ2o7wUw7GeJeUx921AB
1SwN9az6Y0k6u7/rt9h3+jz1kr0YpzWANAjtsNN3+Y2Cp8w6/Mu60OeFrR3GPSSBqPQ630S0jEWJ
2GgQ6cl+ri/+UHpknTcaaE4sggAHaP9iO3eddLGxKgsCtsj+aPiJpZ/NZubjAR1VGiJIiFeQ7QnJ
3gGulUoF461UadZ4w8ScJM9agltVm74C8n3Et4zpgD3NizCIfatqjln8IS/JPnnWGEn4dqlN8kiT
cMUd4fWbzKPop+Kqvrm2DhpVr3eQ7PWBCDBpatTmyqt+xa94Eb6K+wRE8WAuaR6gMQhjRqSdWsNJ
XNtd2aVi8/TVs8ggA8I4bupNsQcjdooOsyccKsnDq6HRjLy8vETZJuQ89CnatFkdk09YkyhJJRmq
JlBO8U1KaW5viyhdbtl2s6pERG4YTBG9y5SELXnuHxrDFzTpcQm+Z48WI3fasCAC+hjghv+joJ3X
QFdb/R/SXOj2JRkVlUfJW73Sf99bzBTuMZn+ySvzC0uXHxTb9i4tu6R2DeCY2c+Xyb2rQuZTc+te
13amQLVDcjbU++JGFHXfV1ZBh7ofFX6ya+IK99k2o5aMm2Iva/l2R7UaIuZStwKj5JYhWuHrFP9j
z18RxpS0EV8FmcsjJEiUCQm6wToxnR6cOwf9Py7Y77Hil3YBngN692zeSwToGUZLNgBz3MEcPjUa
W4+AOS0LN3FW5Zfxy9Hn3JLsBnyRA6DvB6hqAuLYvsqzSyQTrL3srVjqr/6ziIM+16XP3fdR43HP
7CUP8PlcxeXOn3FTxA7k5nFM0jkNItg3Tv635tNMLnEdauAuAs0RTZ+9Bk+7Wru2HcGew/yg/+jH
s6pF/MhKl2uce4jD4khmdJ72TIxtAl5Wca3KyDHDCBsBHZHmE/w5dXLiOKr3IAvcRGquSfDw4CgT
aptSaKo1KQVH2LcaSa8CDl9xRVi0ng+6GDx5TYJ8kXAYr41HWuErXRAIIySgJkTLDoUGnRZstfmx
BjI3JnZyLi2uh0NuvW9jKwf7R3RmqpOwt25m7SCWQkahL/wXwA6FpVBlqLQsN6yFZkCggpRqrxBx
6pXDQ3Qa7K+k4NLyYN1AD+Yq371Vzmfv+tOg61MwWJhXwZebM4gZ0v5uXqQ8hPx8FOOvwlrYhBGU
ewsnniVEVl39/aMURyUBUMGXUKJqWlFgTSsftpLi27vASXGHvP9+zkP3ly4VkFBhsPKEYPbSQk7J
wfD6s0mkrzAT+qRO4uls8d73OEaJI4UuUVJ+9BXzOODUINvn8RODPwfTbLZB1Mdfk7x2AMHqqERr
PqSsUo48/eEdu9/fnzj4Mv2WQm8Up/lG3w9raFBQNE4LQFJvM9gsL5OCZ6s7NUpJcWY84p+pmeYB
oEya/T7UEJh0lZDx1+CUaBYpsfnuz39lxyIqzxN1QrV1fm0hInHfNCdOgp2Y0o+8R7AWic7579Zi
d0Yy3omHA1jX7mK1hnKb8PQCGxNi+q/FsvNyBB1L35GHA3JviSlRqLNbUHPKNQCxOdUPBTaMjtlP
s3hc9MR80tLiB1doWJ75i1GDtIvUXHxxeleXx9pJssesmz9RLy6Z/VvR5sRkuQStRoaMf3R2TX4f
RUbPcpI+2R7lgne1apDbKz3BqswUAF+UEtAeoPYbmto8jx3Ojg1oTkuMYHN2gkfmt3PKsbmmcmvg
6hBegpSDOf8VzdRO6vkPcOcpUbsmVAHUmI+UwyLUQwl4fFzmP3jN/NonselJ3FfGF47vjsBy4GB5
6ir3JqKMInsF7+2Xn2qWzCEhZkQcMhUYqAot8Shio4K89YxWuJ7NXFvTVG9kSl/vkDkh8GcTVgOD
/oEBvf9VZBjLoo0MCaSwSrJSHOqzb/3qdCzDNewM4QPMk5L/m1TJuv7WeYslvtg5v25nVuTJga6O
E2Jt0Tjc95pcqDPK+2hCwKoxRzi373Gw5ETDTHVAPZs8FlXP96qmD/1M4xby4TK2iedLjG/eHn6g
SeIQcVGw9TfZBfcJR7XQvrO2JMKB1lUovSXpfmVbKFXbhIzm7Saa7BJ9nWLacLByPawoX3vpXulk
l0UqsuGabcXOJJ7tsIu4A9fsy0+ZabtVzuLBuPzvTqHXwaxtl7rIBlU2jtU+gMoIZelajtdQP9Uy
qQE+U/s0RwGVrvdWu5bHkXD4s7rhbhFxpX8XlxYcanpwxwSm+Fu4CWTYSyolS2MpLR9dVjDIg++P
xh4/D3at61a4wVWXHNuPwqpIjWKQv4DJPeibEZyDERyzqoxCymPIDA/6GW9H1fOXnr4xZLvk9p0W
YLbakm9212JJnK4AntzzWOCZ1eE5ca6bFzDPREpOKFq/zM1mk42M7RAl00TQGPgtfmMkyvw6d5BX
a2qzUGWNRZoqLMr/IYi4DXcYlew6A/Z/nXK6SUDceQo+vlkssuokIb39V+OsGDK7ZeSRddcevun5
il5ev+LhSQtlpUe1VKFCHZox96P74W9/qtRHNVerfvwkqOeEe/P8Ev3uC7dyWlkpRL3QFmY8eGt7
NEfzeZlbojmu/mJCoAZHqr2xfjUxE4pKDqRrjQ97eS9/dyxZjuQ41pcoikn0qdMoJ93BwMe73bEP
ucsqnajvfgTLeIGYv1ncpVgtgMv3YrbK6euxNsP786PXEhnOThmVsNXCeqtGKGB2TyGHgrqWevxH
gzlTbwklZE1FMEQKb/crioRER7e1Ie5oyRjZNe5NhuMt4u4ATTb7hjgkVnXx3ZhFJhhTfcL5Gg1H
cmlF8NWsJBT1vpSCx8RKCZuAbAu7s3FML51JXI4eKVvb3uyQUggEypn7w8KB6P2osnX1c/6PQRd3
rrPDOOw7/U/tZX7d8J1wb6iMQEZuwECd3qHwqLIZzNkrSgwbLsno5EAGxE0/7taC+tKSoLC7mkYt
NkMd2Bw6fjUOK1M268hvpOSw7ntYqLsuSW4CrfGJvrJTEb41Nw88AAs4wssCa32bV1M8yZpAVPMX
VRuOVN3QBTalCD50P0eUHzyVy5Rz27TRMZy8GRrkKX0Od6Hm1J7lRmrYgajuBeJt3A24nSnncoeg
XBTFAgabuDR3S5G5DCK8Ff7gHckh3D+i6OJ9beXXKqGHyLvPSmOFYJiWleAiCieCfHajIzfgyBpN
+wkw/oPGMt2Grm7e8PzpogwPH02F8NUbsUuxE2AH67ZAKKCHBxRdEGdyztTpEp12MTuCUkFkaeC+
w1zEi1UGOO0SoFm7s0n4ngg88tB7KzXWApaaisXL4VLulY8S21XcYWSwde3KXxMERYtyDAEoeh4h
pS72pXagqwpFgGdqpI35zlc8vqCm9laK4dLx5gsOQN9fhk5D00hHZLraAGhledkNhkidj8JwZ39G
iY45lB45CMG+2NPUzveG0nplBAnKKYvP/YCCZJ8wWtnZPGR1lhGZ3mkJNdV3QU8ghBneWNlQ5bfR
X8zLR1sPVME+S5gcXTGFL/K+s6dtlUZQwPOjqKVlfEM5VSruIM2ik/S8UI5e6xaZ1uLh+mqZ6QJ8
4aK3OjZ8lcscKo4xS8GRo4W2jEAPHbaWBAxI8yUvO3q8BU6Aa2p/N85iVSaYDt2vxshVm7Q0vAdZ
csIkNOvxOv3pJ9aMF9Wrpqr5pGRSyCIXIGGHHNIrcka+WK4PKaE5++rz8h//e3M4SMXsSrXv9XBh
RvAxIx5FA14fUyUAvILG6Mqm5IYn6EIvVzTuydJwt6rlndG6yf8BBKEermRKNv513aGEbfLaMmsp
H70Hz694NH4ATP0kaP1zZhE1ZVTrP2O0pzhpvQRuGmac9n59uR6QPDMlTjl1dF5+DDCixaRmZnvO
ph9G6/aSjq54SaqiXLNDMlyXao/TRPvd1D589PWRmjn25ofpAUwfKfVLsqb9tbofkI0mByueSBQh
kUFjCm/Xa1cZqDxNUjLLjWtfiF4tmLzdR6V+RTan2T/kWFp3FiFYtxQZz9zGaI+P8ILJF+KesKnl
Z8fnTIExm9wq917p0pzItG+8eBEtqcvolCzjYWkykcOfzAfSWuG4IzOMsbCrzori7CoaBWv+T/g4
Lu/EEaGw0Q2njXyXcupqaa5ZCXcqh3z4F3SmKnHVaAa+qX1Cu+SGkWYbgNCNfm91ZS5AzeoC0EaN
kbsGn4xyjQ0uIdKppyVPw/dsSd4abv+V2ceJdt6WD+XMG67QxVPenSQj6d5cTPXRpUZOoCyYPLxF
4nBioqg5Pu9+0mj88U7LKf8X4Y5RvjizbXdHr0b4koLMhKPefilUfiE4fc1S/cFVT+WLg9t5f6pS
5pS1bB8YiOeoICt6sv+U16s1x0O5K8SkPnJQlSCcPqsHsdcw+yXf1i/muOcwDKqbROZGIOdL3xXz
mtQbschxTL57Aej3UcqcX5gasjbv1vPREa8b/4RjdspAQd7XCas4h0Hq8MLu9Hwy2DGDFwdkRBTN
YeBkifFEBLKXaZE2Gkberw/foFxH0nEwga7/WSfMk1WshW69Tj+Hm/6EbrvDNmnE8X8bD7G8nP/U
E4ASTTh9NgoBfoUMpn4Y4jqEuVjecM3dgbzf8veU2l/P1D+dKUlNBqCvFCEIeOUAhwT5DwzAp88v
XAohqjmv2jNYZtEyDez2G6NAeU0qkkgNqYnz/xgd2Q0RZJSkngvZQ+gguoLroPvOPUn05Z+l87rf
Ytwdz9fzXgIe+NEq//iLnh7SCkyQ0+vMV1VgJzdTCiZ6jIkrgYp2Zg/Zo2BxZaq2VwgCkm5fGORS
QeLUhdlTdx2m/vC7StM4biO9vLqAdBADxJn9Ua6QebsGxR5LWYvQveuasFeX/+KMQvcyn7FVwYRK
wIjmVFGaWu6jFIY6Iv60gWXIqPQVaXpi8m+UPxAlxXqL8lVlQvfjX8VwWQgdjETYYWMTczPrHN5q
g/f0iKs7r10wqg48bTTpmkjOhmsEs5//zT4JDLFkLQKVKQs8TW8CmKGp1P3hdSl5KDKGghaNBG3L
5iL3Nhyg4EjNFe91WFSVLIRua04iSLeiX3WDRIUQN9ul+KGaU/ofWNSPlEtk8LpCcHMlpQHHW0wV
a31T1vhdwWVI13DXDVHHMmNOXYqfeiwokXhdAQF2fnHFC40CzD4ZSFwSJRV1NYUgYR5JXeMGdcKn
ijYrl22pCMIDSQQaRy9lCzta+bJ0QudMIjrOAXj0SGnY2KFu9Hf1DkEjQf9gmRVXcHue4BxvQEYy
eZ5GFX3L314vGyicj8FpMjcqeaNbeKq2HVrnjkrBtNDbxZLeZocioJHt9y9iKbw6Cbmh9nDM1WS4
LKIvMZ+7sr5X18EJKBAYeP6UA+FOpElB1zNpCChVpNaeISnuwMvM7ceXBHerFZcfW0gPkRfvrGT5
/4fZS5loNaYsHXq0S8AAQRiyWolgHRPFJ8oayXKjjn3mXNVMTmsQmkbysyI9HmVmnRMXpLShIkcL
ROthfn5QckMYlSkYVPKYE565dxWSbIQF5qrtfmS429TQyqoBMKFOaXkE+Sjg4/ZGw4yCXXrs5wfM
+mhqGxpRudx2eimFxKwyU7XutQ4eUvdyJ6qbYHbeexH546O4ZRBQIfcfVtpP9szRpJ4rr7iznFmf
ahLHgiXnppcmPFtx+/sB60PnL7bWT+JCRy7S9AVWcg+Or38sdzG0QmiKAudZe8vmem0EjXvdE5wD
+tp73DkJN2HNsoD0cKnXQcY5tDyZ+A6/vTLDu8Xd/P+j6qob2SopOiQN4s8vfloJ5vS54S0V2EgU
1KaNGb72pjxRAUfRsuaWq8GxFX1L3lrfTBKWg+q7npKbS20BG6zAleDfXObwkOuFkDl9V9Yu5cHL
MQ4JvXGqE418VPwNEsMk4KTqP7Y9il2VeLkuPl15f+h6zHgjhvXXAEsWi6aJPjHBbgKJpfPyLGpZ
pN7KbHVnT0W0zEjIYjuJrdGOcdlRcsgaT3gKcmGZV2oar4HgvJ0ZDhdQzrgAy1Ng0X17ZfotJFDs
yrNoelHncGrACrd7D8TkPYfabQdSaBoQmynvi8fn+IjUVzT9Ro7MQR5ip4bdrNjbUTEZhDAfl+JA
hfMO0Y7IsfRQlNFM1lO+hw1Has59j/rBP6DmIK2ScInGqN0UWW4kkx9+sX82XLkSh47ocAYWDAr2
KLfAEDT2kHDawFjrRimJpOzCpI6128+Ro+/UhowYFn9FivqZ3ph5CIhQf0yYttwod7c6yFme/zXO
nCC92jDVaFsHfdRQFhDQ+OveUbC5yyojGcPHHkw2ZMuzH5qdTUOSimMboTd1DK+6S/4C/ubcL1FQ
R5LK6PmF+3bm8fPIFk5JOArti01IU7BrS+R9vU7d0qg55lvHOJw6ZvVbMIvWKc6WOtXOos125gxY
0vFgXUjxVw+ZWGh68T9Znh+PSVccWDWJ5iq6atG1aM/+EBIFsgM32Pkp8z/BkYP9XPnGj5O2VAqS
r3AgIKku7s2SLuBJe4OUWSOvv43inCBv43CvSbGEQPajUgKj8+1C6TjCQhzcL/9bnWwOshQgrb1n
tJYItzUuniljun/+9c9dnbEH0Bu7keDO4X/9uOhrrL67jQAWpZle6mCV0YkIuKtDeaRfMgl4pyBL
riGzZ/iDrMLl0/sNcfL/L9WPqI13bVIInXdThPG0S654QxowoMIGPtnafFHSqxT+kGaqclSOiPNP
cb3MTcCNtH8uhIakFLWx3xFd5LMNX5eoCKY5XLEdQyDxqIF4WW7m25KC1CYduhGRwg5y0M36MpWX
aLP48/zOnv4SklTntCv6Xk4KwMkGJ68EVKiGDwTmMQuKRfBuI4RfHUrT1MLRj0bpZtb/BPt0hlbB
nAyG9YiDf5/j9swSb6Y6KxQxbrpdDjWSxRzDiTq+ZHl9pGbiMV8pvFESwxlhifnpylrjuIeiUvCt
RcK9K94gTrl9pVCUuRIfDqf6/oxyRDkwSkrf9GehePQ3T8LHtrCagzKH42rASE4wp9T8EEbXDAPh
tvfZzaf0wDL7PM7k9i8Jx6HD1M70CJItcepiEAEfMGdE5coOfr0lh5l8A+HIJwQU6YdEMybk5IJT
di/pvp7O4L2F1Zfv5WW6mSzERbtTxij6ngM3un/HTf7yWyD0uzGFBCLYTguRX3X6iR1unEp0cROU
cF4QC1hvVBHJzDGAIiYwoQ1QA/R+KoXgMH6oPwsM+piiEe3fxOX3kllGE79w5p2E76/V1iHdNvGw
J4VKaDYLR6mSGAbvSkhyIEW6qInFiKNfWddzywEhDejacz9TV4NaFba3Balyp08vNW5dh+y31gc4
T9ac9fvJb7asupWFukOpf6sDnzCkbyEGRqrfn0n/y+jE1KtJpukwt/N+xvsWS8kLhzKOrUIU/qeK
PugHQ/ROBhDph2pcJyr24dvA57GscVZ+/iGSbS0Yg7WG4E0cJSHikQoZCFS9iXRlkefYedMvZ12y
tJQ4kca3BtUd1b+p52WqQD3rMlRZ6QMGokpeXY9PLf11746helhbRAhfMmcH9JUBZ6rGqFFam1JG
XJl1GbHwikd61vhC6weYbdjmbakOEgW2s8xoRP3BblML6cX35VEYJVthOM4fIZFxziImE827vQZO
psGMTEmsD6hX3m+rBHU7cOMWoX93MFezDRJG32IAnZzTH53wbleND3wlJcHNJnPb5pIrhZIa6Ojw
ogUzZ85BcYj2oIuvBidMC/d80668GTQocHlgFh808GOeSBO/FuzvMBrHVKy00eskeJ/K3VLHuik7
9VkIk35OduHC6gJuqJ1/y1yfc9of5w1jKGYfEsuvFrcEO/CDHNOvR41rIivC0oPw8u12iaw+hWYS
TvQt2EDkXlVAYCjRccNCB26+jZff43xAWdsiFiiy7XHm0ovhGUHnAB9CRFO874Yi5kdGtIdCTHSo
yi+riifxQnIoppJMAAuLCBqPbdgED+7uvhMm4+p6KnFC8+SJzLkS0+UZoenePy7lKiWuKmcUBYEi
9sPEsqr7wh60OOsPnbwKyx1B9wcMjeXyPh61IHDJX51Hubkxxp37ziZ/6aIYO5o9/pUTmFQoRvY/
rbqbMh6O28Jw/M2F+yBgVHW+joHEXi88lcROtcSjQ1e07WEcYI0IUNyQ58Tf/W3yf5lELYraE2kN
AEtpi1MLS/E/KYiXEB7Lh7SOZaho9u+d59aG9A5myIoLl/DlWBLxcbbv9an4eMhXCsnSzpSIGv74
D4fN8phI/skfIdcIGUWWBr7y6OoQKwdpLmtRes296CdNUJkEt7AWxeIUvXHIL6MvMGJcioTh0PF3
MJiJVgwbS+qJDhykQGoudLcWu+xc7r4Gcdp0FGNDw/0ifgsSDocE//xEeV+F/up72Xpf8ntYY6rO
ZYeOsBayMKEF+gXzJTjHwBxuRepgJBV2toszVKNmzd6OOFvsMxjAUlvDdI1OWjk4lME9X8v0VwhC
4EQ25ilDXxh92gqZ5HOhkPYBPD97uW3K618lCQocdRKAgkkqwvUU4+d2BnhPZP2DWtkVVJjjB7Oy
5vW+P5WH/1M8xKCJqaXKLoA/eqaNTpvb2Cf5BY9NrWUk0iG7WLCa53DYkvmVvoUxGSzAc7b3jOfy
E5kGb+jA1ws8CuWCSw4E0XAUZzTq2iTsgjXamGFA8gKafVItGfz08EmIjcGRfKp0pju81/dpraM+
hAcwYfaVfxcAqFTyh00w1gumB7Y5+unnJNEJWfBVMheD1o3aX65RnUgEY2pqYTAFdmPmhhA29MjU
5oyFKs+Dc4+Hhy4EAI9KkTjWQNHJR74V74ZStzmAPuaQSrfokeHTbUhKxDoMvwK+HjWN/abJHhNH
rutenifXeXoiQH0OoHuk9qvcxNzHPSe7ULhi7vjplb9lsMniZKBoxHTMOjV9mmqTEqKh8GUoOJkn
F/4unuAYQ7kIztYS5cNEL2uCDBNoPNp37vSiDL2KmXIWJVlQCO/TxTO/u12OR5NBlnfp/J0SlSJ8
Oo1xfJqpcm4zph5tgVY8WeQGQOLiWtxmZduD1gMRRlp/E2Qim/pesC4vRlwRhDj/EPw0mwCcBq1h
lLkkKaK+TYgtsKnyTzHaQCuTmbSMEzJl3ibPe6XtN+BM/OUskOqw6o1vclaUwCrmf/iyAjedXnFw
MgjVZQqUpiykX23ArcTr5FXHviQToWvCpjhUaZT0/ahjc7AiMWjnQf2dBP6vfEkbtfKdSMnJNESQ
2nDOKIcn79n9oE1IwM2frWOaA5JrwGtBnSFl7sCFVZ8z3cXp9YBQBE7onZcpfHZgxoqscMKltVfa
OZoGGvD8ph3SPfpZfEhq2L+lE0nP2i9qH0IcchP1DjOv86E80Yu4CGBaANAjwjRpySSaKE9BKUg3
rMs1JYoZNcjzsLDTxGsvKIUeyggDxhQhpHwqpdW1YXv7UIOXyhN/y4xkwQJxPmreM9DMGLrAtfTm
7dH+V5ycqKyfwWs2z3MU5CHrc9qslY5EwTmQl3M1KMqauEpsyOD9zZlXaAgqIdyynacXM2G+xxAB
4qAmGDlJijStabZ6ZyYssBlmahrw2NMlqGO9GectZolk+H72cs4xIV8E22waNnzDzoFh9UPgsQ3V
343DqfolpXlypXYpwCop1YH9OVnMwdxvMTdfJnTA6PLGhGxkN3KSKAA3s7AbnX9q8HIwH4uwSjxC
dSOAkFUcDUD7Rn9YZbZDTWRGYhCqtJVvEopEzFwPMATU0un0yIr87WXGsgzgbq/A+iWTl2yV0lGE
umEtVkrBpV3qrC0OTobMm+woX72MXKrxZKEHhAKDohM1W1mvH6cou+phc6N5+7IY0Nu+xozl4Loy
4OCdnx3MMXl6b2jG8JJRhBc3T27SojLyZonhPlbtcWw++bUHShfJcuXhXntCBRUa8UqrZe4mybWc
VVJRtHo9AH7J+Qngbhoqt7gN2MdQ/x3B3Xjjs23ly6YD+tOEhSYj0f5+y5hV6cnKWMCm+shQu/uC
TqyMjT8vwWMV6kPbnIXg8dEdgd7l1Vd6Q8XhBjzxyEgfeWiqPHKODP8zUsZSYSbNqlyhwUp2/YJe
mC69R+YtGeXZmq3pCdC4bL83jI3yZqCthXccwBQnx0MjV4ghgbduIs8iwIz6UTuiYR2Lrds3/PmR
iztvCjrY6WxyP4Y49ecsqM//28Pd0XZgtv2pRv1UEzyZ7ddoM8luwv4L3ArTZZn/r9SqV++5EQ/A
0iF+pFSeP/L9vZ644eFxt5c4Twku+/elTFzXf7BMCleDLqJ34J3jMXvxpunKY+E4QOHJ8JaeUcEh
ulvKjOTW5ebXjKsGdVxVn1xf9iVbhwsCJrZyWcsTrFOmtOnf5DHM4C00ifpkME28qZyMje2HezaE
flJo8Nt7M/wCKTsjnCWoYPFqKDkUfFtcdox39LkNJUSwQv5mHJRo6nXRICjLuiByBqxnmMVg6TBG
kUxuORFSc9/GuEjd9OhmaB4zzVzDSPPLTSsLvtebBfGBQiutIDwDeevkyqOXQrV0ZFmrohwgvWBc
ATcm3b2JxXjpFrn1mvKOPOLzYvh8XAqEO71skiSFHXrHoaXYP7zXd72aPlaR8n6jsH8KliBXEMc6
YOFPrcfYM3Zm0sCW/vNzmydhCp27zU7NBAAQIQ9KMrUFJ8hzdEIyLC74FB9kUO4oj7c4xbWsbWPM
osMLgMIgZegfodc2E0KzTl8liO+1dEArTAPsGpONmr0Sa6p8Fc6K2W4Rr4J5ckzC7nKfCOMtPlyO
6IlwV+XFYMFamVIqpX3BUTdx9DHss3Iu4MhM6RpO2OYnrs+vIqmBCVWds4lvEFd2eRvOQx8I75vJ
8JG6Fzi5VPJ0I2CkJz4OsUcjqAqC4I9TueLx/Anc/gr0Z1dT/M8Q43vxbsNwcl6sSktPZXOHDC/D
FYs017b+KjAWYEoNHnrgGgyac9OQx5rtaKxzWe44JpzvK71L2ZMyN+eKdeBOwgDSLEV2gdJRI/bH
N75nPrGa2JaISXJJRv5qCyNUGLGSYdSX0FOL8LQ7pMK4YKmectl638iwKDgidJj0bdsP5t3M7fRk
Hn5cLZAnU1K2oKQv5bm4pgrF9voRpJWO7or6ZPJyFfSX2mO5Z6xpDRujX4ASivPO3+ONLJYFZc9m
hiHub6LmWKlWVbvYOtNRRKu1h9LaZOUORtUkL/lDVY4PUnNsotvOa1SPe4ZpWgv8RtpKFZfI3PBq
atRk+8dysebAIEjwtXPSu69QjiJhCihwehFGLsiZ9R3fNk8vESLSQWfSmCQglbsTpIEvGGupf7GY
QNixewvtow/QkkyxkeMsDKfkxdDDoKO5wWM2ToM2Sppy5Sg0wFV4qqvoR4MbDHn4Qb7CG0iTwztv
S0vuzaRMiUOU01VzNScUR9BEwNX4pUd5PcR0u45SDIEcS16OvsCnhlH8i9a22ZyXR0uFFxc2RouS
lneo53tGW/rhEmiK0QfzfpEZyQBYc5vYhY3crH9jNgJZtahW5OXpoYYtnB+gX3waBOzhf4B81r05
lA0hDjfHtvOoeQgGvEL3lNjkWcLFi8+xoirvsd0RlH5pQXXrQtsL6/VB7GpSZzQ9M8djs12O8xiD
ab/MRSsspGTjYVAVL9riZLR91rUbuM3sSVErDKwQwbLGka80ogy8zDNTUsHIm4b94iIjruKjIscH
f4h4urGrUjhJEaFiY6TG6BEc881Dum3CHjOx1DxQJmEYtXSJpD4LBPXivz0ml4uGI9IkzmLb4ZkU
YRAaQk8Zr3S8N6TuWg40yvUmcEuvFgt8Omick1QuRrGKaXSP8L0FNdaDeZQrqvdawJUaDar06BIf
cuoakYUGTomRizOancrof/lCpH0JGwONSBF+GQ9CfvNS2PS8cRH3VT/4hpf+tQqkyCfO5ySs5pd9
1laSELHhY1OsZOZdjOP1gTHJvdSg0d6yju5A0EUxHFEzRgTVJ5NTX2b24xYnvkOtlgsQuxGe7cd1
JFzjiDIOhP3YuQbzhaPRVxS/DXaXC2e8fog8ly8boSPHaku5m1WGbTil8SbzWrhw9fubg0wKeyJj
CABuIbXcfoQf0gfn/+nZRLHe4J2JUDI48Euw6huSW8H0Z+DnOGbML64pWTzywywnsluxX5GgnVlT
hvmQcdFdY2hytQqm7iIWTYd3auhRyfA1rCYSYHeXnke/AInsTntR30Cp+Aj+oDVJ5pFmIAUFJhPF
dmHOe16k0kZQxu9eodxoQOGUOL4rKDQyn0UVGdkQYobqL3Rl/pGE4zNYL/1HWXqtIABFS/J9wEQC
LexXdCJlswo1+g0VBJnusOr78CmaN3+M1pSBOXSmwXoBUSCn0eZtbMcsNdzBruEg2fcdb08i5/Sj
xzE9NYbo7ij98F/WcRSg5LoAVeHOlDk8e32E4X2Vg3mvoWiWxZLtnIxuuIlrtU4VtitdhqtdVlPK
KjyiUgvmsg9TS27bhBeJnJ7Tw9U+0apFJBGBiThfg4eLYBglMzmPJT0a7PLo26WNwaCfYJUxFNCG
ABEYF4eUfUyDhNQIYDNHhi+PlJk5ZP69iNuW2Sb4xk/DsHQyE0gBjgMBxPq7/bKro1lhYNuCWGmY
rF5KFgGlpL+Za/iO3mBy22+DwppKEDXVK26608ZEgn0+DlaLDpPM7RAARYghJmkccoYx49fSVOU2
KELz1T0Sqo0RxGcXLoyt88c3wBlTRuEHDM+8Aq9x1fQznNF5S/NP2413wWmIuGiR9NkwQpEG04b+
I4KJ+1qZQX3jvhJZv0FByiB7At9VUXbhy1dwKaEXugVsekeEzpOL8FyKX9kmKM+f8WEgQs/3Wo3X
hxFIvqASSalWF21A5QhLj5gkKk9irOEPZYii2reVxMBHegBdp1Wkap9/lqHNhX6dIPIWhLdImheZ
oW9T09ZKawIqVsey6FdsSLlkeBlNkxlfiloUm3bhPOB2SkflzxdV4GFmxW11eMasoU8IO+mtowBF
p6EZ9C4lFvxXdHwunh33fGnj+7RtMkW5S3ugdStPiH6faM94Zw04wiErT/EhdShHpZSlHIN98qwe
s1bkzeO0O3YPbFU9Hq7HnbizwQ88Iv+ckFPkbrZhTan0D3BpW0mLXJWxDFa9m5v9Vah9vgZTP8+C
dadjcQ65nWqnL1Gm5t6V0dR+LFMQKXbfrB+wQ1zTLrYWIj+CDlO6zePl7kREgLjvZQgeNrzqPAkZ
Y6C2i0ADXOvh3ZF0gu6Ioz1SVTdXNT254ayVTw97XIPPc2N3S6HKE8jWLDdKg3IBo/m0K+u6ocHO
EfpN3su46H4RKeDvhSpBYMhBnOmHtRJ1x/iXQ/gXd8s81o+OY9CYz3Iz+JsdaKfXbezEKAg+yspH
3FzjWGTEYbbswi1xw0TIvkQ0F257Gd6UJ3Z8gmDE+0BMrjmaFiLIGgiHkaP8d4uj+4WZI3xLf4wU
LyOWY1YfB1SIl1XqdJYXG7YHsNECm+/4GP8Klmz8ZLtPjNvfuDukhsaH7OJGF49Q0Z5jq59dTNdo
ksbFFhynveMyq3tGh2y1p5WyisocEua0JAVc6MTdYFa9g6E0u5NUpb+OdFQ3gVc/wi4o8q8yPg3K
LJkuTySBscIoD1FrM6TGDXcrQzjjwmwDI1MHMBFBQnfE+hc3MNLN3jEV5Q2QPbrSTF4wFFCSChag
gYcDpj4flss+4HlKYEenon1l7DAUj8jATn6poGw55bZ79sKUY6LklilfTO80KjnkdszJjBvv6/cn
jrAp5SJSLJsWiE3K04Oys/5OeK7VO3h3PJleCPzzh242ScJA8F/V2CNK0rKgY9Y6V8GWfpcKff8g
0CyL4vYHh61mSFJsCK98EbYhAR84/awOK5hi2+sPf9chvaU2qDw1BrXGx/ay0BBpEJy8dxUWMhDn
s+8/OKQnnkFBdX2E1BoD2Mm6BHEZiY17ZxVzqtDRuyt5e/2EfzF9rELX1NDZI5p09jTgmyJfVqPt
USezYrce4ar6rLlCRmFgVrN2+J0ZzLiqGJdIzkYeZJyamVdCsp4UK+zMf44y/TA1+klRjw93IRDT
YbrSXf+b0RzDX4HZyuAULAUCMb6ZJ6nUulN9qC1XrkU4k3wpD5axNrJpS9sego+AlHGajozmoi8J
U7kwPdcxZuKyIhTZONzFz1pgcC3VYuQL+Fw3402q2XZfByxtKvDb39Iq3KqTRGAhnXkaJxWPt4qR
cSvRX5gZtSGsUTDYHIlkVccLq/QaADuIlCQuwXd7AEz6hunYIzh7Njg93huAgPlqq2kxQ43U7Tyv
H5qnFJ7zTY+fpKRRarGFDMASmU4aFis/uqepPu9IzIwl38ZLVBEwYrdEmqsP7ddwE01xhk2rIZwq
gAHyprJYG17t1FiW0JLeBaswsTBIzTb6Vv0kn/QzFQzVCCdjf7MNRAgjGRmLEoKm66NgokTudcvz
uaIT1qbZKcvUxUnmjOA9G7FKxp0rIMg1TwHs+Sa8fIgfufUKt+YQ+2ZP3VnGflhRluYcJkxeYI+w
YoWMQRuo6rVw1tf/RnjOjDi6xt7oCqUu5e+xmINqNGg4y1IUxKcN4eY75ORKZRq2UMkHOgsHcQoe
awQEU85p1bqOKSGtdOELfCPLJENiZWVnwyX68N86WbW1Q/s/Id9AbQysQcrIRb+JaJvXVVe358cF
TjEssfY/R3z83MvEVXYLVp+5SR5/q+rRZZk/msMoYZgOqJRxW1HGEtYmMx4+pQuvGdoO1fKv/BvA
XtQvi2jvSiu+NTBkpxHEVFcxkU5fv00hNKCBlxUXLgUFlK7zkSjakKKtEGVTF7heqh6wqmh7dklR
k89BquLJf4rHW0PjC/q9E8tSmZU2RcLn/z6VS35gdEreJjKkt0nE7BD7ISU8DagJZFXleMBZnNyf
jgW5umVtySZoohSsBRfRMqfZs6FUF4acT78zLDof90eMNAiZdUZIa+5Y0NRwAT8vpPvFcat+IZAQ
MEBvqaJt72pVv9HebYaBnhi/8iORLdd44d2jELiQ/XqwskthUdG8ez94B2gtqE0eEofW8YV8T2dA
iz4+K2ijBtKb1jlJzJr9VyDKW44ogAok3obNnHHZlINktYPnKl2towiV0apDWFxO1vZ9fVevA/xL
AooRerQE/pJ10X0Egj7tcq0rf5LUWMahrw11AnoeFagXYnSBrYW3/uUU0FHio2w/GFTBrZ+oQ2DJ
wtGK4gpRVL+VnLUFo0i53es2t7LwC0d0aeKBD9FZAi9X+ed3MUduinz/Gu/mp/MrA4xcB38xvfVS
yfQ15aCKf3HELplZrrXxWA5l8zOjonZ0g7KXLTJvnKv7tI9FI1l/Kb1/fGdzAiec3/2enLepVB12
rTpVHZLcQJoor91os+t4mv3ML3KNtMu9HOwW12nZxP6HDvLAkTIn/X5ydiMMCKYyoMwBrnYd7uMN
XtgSG0a8g4xM3Tj8nYltFthhF48Scr0Yq72Se6x22COlsEFAcgTdng9fGi9oLzGb6EPkpha9m9P4
R/VkrB59ZIZQqH5DwwFIrCGqjGg4fjfBdqdey/niFd1H1VlfRsRfbiv3sB9d4zWEo3GwMj5GmOZ3
QifzLEEomcIHwUBT6Pl/bkb8gy3nfbp67xp7+o+Dut6z5bLxMWPyFde/6JMMd6yYX3hp5RrhYMRS
Ev9hfGuoTQCUbS4ETlfm01suk2n5S9vCE9wkEPG58fblduIa+hRipekah0u6n66qZzQ5Frz8X7kh
ekket4r+LkBWxZ928xGrIcsD7gd1vAIbjVoOyQVLQh82x1PNUZOZUrnZbDFsE0scWzDXnrgnH3q0
X6l/oIYf4pKeXsjwUmGyKu8W/rLvQCu8j691Ol/m5DEkzSeIr3RH5FW3gWzV1iwFjhUqTACGIhIk
DlbmcsjKsGYRRK1f/ZnJ/CMQVJpLkKeZbuXgpw1NOSFfhrSbW892X//b8zsp8s/eMddnuy4GoUyH
DphGpWOFH0/TuP+5haLex3cvenaJWW2uDG8TqkwNV6uvcujTCNvHKEnGsx+FlEm8Jl68lb7K+cHk
jerNEXUG/knSStQHqio5YmN2AKawc23eP00K93ssxuNkP5xfpyy1zKqyOhtPW5tyqUNHk4A3tlFu
aFMm0+S9o/Bl8qUi/w8kdHrQm+jUUVH60lf3BJopgjhZ7xHPLQw3xBmZpKPeqnK+q0KXcrLrlCS5
hrmJBHtHUM+enTJO7AMPB38B9ft4nY63/vv7IqMGF9Afx3kcfA7E7YodO+mvtUd3WOLmSPWRXAsB
6QHivT+CSvc2s1Q47gOJ7YnhUXkESBpxDRDzebPHapVRVl6CLH2mw+gyINPauDEgSUsN+dr7cIO0
gmOojx3E0c+Z/u8SpqGYyM5hFOBIEa7ubak6pNX6Cg7rfE+Na9p9xKxP4NwLxxGv79udVpZl/v1h
DiERQG7sx+Nz2qBtCe3bcnkRXCdfmsrXPds0zkmeA+8iTXiKs5IHgHIsmqfggtLTZv1C6/xKkw+O
JXPyjE/sWmyK4xQTbi365dMIhPH2llJARWIlcuJWtYVh8NjWgBkwzUL0WFB9kwQj5+Pa6P+UmUJy
uXIumHUsrZjENGtK0sfyTUn9xjNGNKvxaxU9eKKPyzZTB5HDg1FBAyDyYdnWwE4Q1LRwYbHINcTQ
zyIsca7QixAcTJZ2VagahQehMn0j3Q1Ka4x7S0cs4u1lAtg4zEL8eFn9/RIUoq77NAXPae2WjT48
yqnlummV0ZuqlFVdGbmh+0eI1DgPlA1w40YXVsJ1gWXyebHfX+v6/HEF9puR+qkr10hF/9IToibZ
hPytBWridjPaPyTHwevmi0fjll1xdRT0lwwsbGEX+/XmkdEN1CxqEpkLXhwZfc3kuWyDPujg1Qzb
bKOgAukmBKQAK8+lxTQsahfOlY7Kq65iHvPGs6kA0FFFp6YyMdNGn75/d/rw82We8GDgCJJO0xEP
79PTo3E70aSwlJIQ67T+buDYtd75ZeoYabRhgjvGKI+jAUL0L2ndox0MtFV3LCrWSbhwqErWlHts
w6gZNUU/L38XIVeKw1rEcVRmGrqhuBtImDX8vV23qA+cKI9LIn5sr3baNdI4qn8Q5BB6WaR3SiEU
xIjwDkDNAHgY1H2BoC225f9Bcerg9qt0UYwadk5lODJhFN/Be6Kt+wiX4wgcvtF9dfue4iaObRdM
QPquGUeXVycw/z/p9OOhi2m2nhKAn+IZT9azdqADEpIY18nfhmNrsolXjZBUJeC4WHva9gyclPid
DXI+ckRHKExpqlFEDz53qUv7Ec8IMuPewxC8n1Sqp20ruvjgeuHz8u1E77NZPjQC47IqlAbP6Qf1
yQvnWphwyTR1WwzHzm8WgOm4Ruju1P7J/iOdxIac11ahutiffu8VE09dCfQFPNQf1IdV/aF/yM25
6xLm6MMoid62N3u5+hEJq09D/L6AGxvRDH8sd3OyomqIu6EcI5MqDEuvBWn8LCLD8aWMVrGuecjC
0sQG+1RK5xzg/50yUMdbG2qvmuAiD9HYV+i9JPQXdrRBCUZgaFOX/ZNZfmNm82UpBZRgkEHEkjs9
2sc7g72uxaUyyWMhFes/CtmT/MTa/5X37bE9t59+lGBHK2rgZOZbyVmm0SxkUYL060bcLjtykrxk
VgmDkdYtEj7YKldtjV12nopT0DF3mLWNlxe+kkbwx1M8nXEF7lbSXhHyFxFTDhuN9j1WFhcgaM37
oEwL/kJ7KPGuujCSTR0hZsc22b4LIT7n4MmUYj4f3Od44utmySNiW1AmK5km1NMlrPWG191HzwsG
I2yF2WSFudKahWtiVrocCUvYPvBESC9T3Cs+MCEyfPZRI3jDrudsQedzOPIfW6qoOtN4Hi75boVa
CUT8AP87dxaAq7WwLgxBnEwVSIDWdEs+EOAFILlB5lEBk3VHoScumqMJRQJrtIpj62e9S6D6VBUs
sAIh3V+8giBo3dbXnpx9bgMNSskesAOMVQmihXA4jMHpBBeyrY6A1X+UyCcnr55+V6Rf7xYt5k0G
ZyDlCofJa7mEriClfKvK0cYPThtT6Rw9jTlLd+GoRbvpoNnFkCWB55a6zUAQBdX2xq2zUtmb+ujA
8wE+xoaAIl+JSJb00DBZ9EVHud+iaaLHDnJoMX2LqfxMWLCesaDG/SNJLKVQapXY6M6qnhnEB6hM
WXDIYPMicynqazBmTUBD+gEEZrqEHoDkSO5cn6WZghn6lrd1fbzgO5nbnewsZZclEuzRJhRAOTo0
FCORz5Kg6Ul1Ynlpd/A/sVHWlEQnjw7J51DvUA/KnQhoBYu6Sq2KmRD5mKS0jKiYdIyYSA6MmPRn
BFctqk5wVvx7C8zJwxGXeUo/NZdS+c3CwAIKodr8BugPJwQaa7KM9AJBUVSUskZ3ERAo43Lc6HCe
N2QAwjuphtysjbki8IFLUA18JxPXZW5ubDVBMHpoLMEAXkRLbufRltTaCS/2xsrdKeFcFHuWsAUg
Mg1bZRIVU28Dkpi/LHm4stI/o+mabJ7L25iXP9JfTYmSTgjia7DGERc+5QMlZ6p4N/iW9bPxLchN
VOqTGAr3wCaScDWuujMsVWbVXFBYP+amQWKqixkEmnWHQ3tnh0OXOg0Q44HQmwaeEevSwgGlFiFb
lC+p8F0g0FX0X7gvsR46ga1GAyRTCUzCgkwxp2tgdbUzeimBXJiC+5gLisZUim7/4dB1vwGbk6y8
CdmXmbPT+1RKbZtW/GeTUfvEdNffetL2QNMOlshs71P2QBxxZ0Alg79OfgJQ2l69L14ZDgqKl+us
2HTHUTm2m3HUXEV4PsLmjRrpu9WgTNjQQw2glPBSJ7S2z4emufwOhw8VDByinDdqFIJCAnDBRqqK
jQwLJV0ji/0Xxz7/D5lvfEtmv6Di0CqTTcNIiiIJsRYdxWrY2cdnM04NohoHzdIzojWWj4Kfend/
yynJbuqE7Y2EHo8R+OKQyh/Be+GfsJSFXxGI4Bdp+CSPv5bg1SBY4EbhsgF5gOsZOKvJoWDSY1ne
7DBwXchUsX3ZO+MSfEU5s48+poHz6L1nSnqQHoPFMlYdp50wmxn5mldhDJ7GB+hQhMm6exeDEfbh
ecwm1MxBaKejRBZ+QDqK2ZyCa+YM5yE+E0ez/8TsH4JaZi8CnBJoVDl0qwPr8YwrxQ9kDDq0IX3M
TaPMPwG1lqUNomk+E51dEeeNFmlRr9e0r6U7qqq7lWrUIQ3gWpa/6SYdZskFbCaCa0kcAbb4kBaB
StcdP/6G8h8RhoT8jiq0OCteELEIl1B2Xs4dKhJMo++5J9djtWGIoMXPzZ6NVwoI4Q9E4jwRphVk
iK8fVa3SWrt/tqDamL4hrGWxMoMUGqsdSQW9Oqdxj1Dd2Hh42FmN9m2oXVyyjrWVQZsxRtG94aQ6
O1kskczfDVb1Jph/jk3uTo9Yp5z+Ebs0axe9otx0s3ICxft5Et/ngzO2u2/HDuo8yrZ0pvpei2NA
EXAcCEGiT43u8+Cr+u/LxBgcYTMGFMehbExcaW62PFpSBPz5/nGPe/ZQbW3ics1Urs3H/yr8nnXo
8oHQIgFVPsNZTst2CwQJ2DCvBe6cABfoD6EZzIP18pqhM57nui33PZ61lAWbyVLeMfdlf3aZRHgZ
tEbkBvNyMfY4DEtbezxHjrtyr91AXP8cUuTm8DRZZEmiZ943IZc0XDUC7Zhkm2cROsdlNRkXyPYs
zH1Mog2s8THZu/nGOQLUj8tTzcmeTbKOakeCzImgwYXXxktuJBZaHn9y2ZjalUl8CoBWkzaHEgke
NK/TIpeUWhwtokj3gFN+Ym2JE0nuz5XIzyAEtZLlNS8kyU/2RzyoyN4vKJqFBwwAUp/oH3DN9Je0
DGmonO7eln47KG3Z2iHRkqvCgFMgSAPyUzhH38o8qfoDpLbAyCqGEjMyqNU5T+lNWoW+QaxWq7iX
U8n8hKAIht9i4N/WP+RZ937zSmR+VVCy1LDl936DwmlCrwqEHdiIjafE9AF14dpaP5XzFN43SDgk
oabnMc7iUAAaaOZLcMRh8JgSw/2LxS1zfIQ1XGkHaAUvRmYd6+9Q6jUyin3IlYLZLhidHt2zmUw5
iAt61AORhhFC+0n06lFSMNBpoYSQOpnKsnCc/vcP+WHYtpuqpylOimmMVYRB4VtKnbqjuK3QXg==
`pragma protect end_protected
