`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rQVIWUnVYlNYBBRywq6Mr/zlwEmXXvqosKu0jSSTWIup/YSsIfvrAurO3yl6F0fg
GNmEeTcDdmmMFJDypHAl5pdAJ/GQgd0noorAqEhC8N5GROYO6ACLjm24u8pD27oF
mWJsvzVu8Tkub/d2HuJ3T7e8KTxNkZhiwMT3kOLo18w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2240)
LL6rhjPg5IOzlfp+htySHAZE6xfMv0oKbk+6Arwcph6eapGBkgmFsZmDs6hRBMl9
HYo/lbj5RdMz65xUtxS4CIyvj8kHgXN0XIfwopEuuc2en1K3jlx0ig4NT7GsFuuo
kVR8oC2+ePQZm+XNTfFVoCqo2UEdK0XPYFsaGYuwvUmY3TQ3wQfCKd2GAVuFoaTx
HZvC8nyIs/ZPP170AkEcRjDjMHfFMzwz4kZWb8S0pEg5Fc5IpSXn7YUUwfvzwQne
ZvMbq1jdk9U3aGFuOgeNvuvuqj2S3HeAazrTSZ9WHOF6bdcN3GJn2F93ouYNt5yy
QCWCIQexwB+ptX4SiyHQFrlcXrJKL/0zukC2qU1nQzi0Ahmp+HMociqvDgszZxP/
w7ZbTOhpCTGX8Y5LlqRyRGzp2arIZigG8p/mNROsRJvlZWs4zBiydG+EL2jCSL8g
+yaVf3/35EaLgzkNhzevxDvhxIHM/zQWgXPCnRgiikvZq/IlAxlGzJl4QkUN8xHn
myZByjmhGNbOWzS9f+hxjoskwdTAxkXlZy96J1rwSxTlvollhPKLIfyWaoctvDSd
ZeO7aAAnR0otF3t37zCIzNluH1gb8uAszdIZVrzGklKubpwhgPTByLJUFd4aRFsT
5o8kdFGlmOUj9UcjGBfNoWHH08VWF1v295bVKcjOzjTtRUWiYtikkx+Jq//6r1fa
PTB1iG7v570eadO6apHTxI9/6USCH4SXJvh3HJ9LiRoZJnygx5u+rtS31KoJvM5O
6T0VLw0lKu0+oPQLK8LTT6Qhe+d/Gvd/UyMW8/kxoPNOiuO9fcUDkh8sm/wpV1pZ
b1WDjAHe4CFo9gZoqE1w6ODSBaPjo4S/PZMJNSXl6eP7J2ngxyb2UeThRZ/B+D1r
t/gfmkqmT2UUPsVqF2y69uZ0a5MY5+DsKHLiNhCyxDatwcbeFkcb936cVj/8tL1P
93SF7HnXmJPQ+lWxxywzQuMeFxmxRrmcIF1p79fbWKg97wDsFLSblVXui9t25kLI
3mYs040Q0eEYiyiVWtIzfT30/vxcl6mYypqeuhJIkHoTX7Jp4cVBZ0gOmp1HuHuu
FaMtekzBnvZ4AzGAY/FWb3HBZu78CznNdOjLpmWeAtUphBR8VFhasU1XDOAQi5Jx
PG1egwzZ//QOEL6/QXTBkzeYJzDXQMh7MAw37v+AQ6QG27Li7+pbneOAlImvQn2V
wOgUkjaNVkdvxWHb1xDzCm9GCBHkgt+spoTvlJvDmQ1A7IEc+csaXdNnfYxHGlxt
aJp+nL1pVf73y+R+TwzVyEl+4XSNWQFXbOk6sYw4vQvO79r0q9ifn++ltoLi96DA
tnDKvd87RFfr1WRDg6NaJad1mddt8GBvujYnmi3+oGji3YApzHCVTLr7fZSDXiMt
sELpAzYFGuAE2cKM9vac98ciWXCVlJNR8YnMEsz1z/TEJz+b+UFbE/D/DnWgUm6v
Ag8gN9CIJNFgcbdUekG3snMJnJHX/3qDWpY/nA1TJBiT+Cu5DYg7fkuA4gFSjJcb
fymlQR1Od/F5/MmIDyHMxg/BekpLbVTmQxs+/WPl/PG2bl6ALDU6808cCILUCVMS
jhudqDNLEJ7AbgJfDTLibkNNoBmB7vsqyD1hht+JqZyzfBCI62j0gYPN8U3RTngN
RlK8IvI0KwOrlT+gomCMUdARyF5jSN7P3BcdvBSCjHAiDx784AcK64btihi8DmzU
ntpNGUWpr3IX5BEsIefA4/9FI9/erLQkIqcUkS72mPbsH6dhjXg3MvZSQV2UY2AZ
X3uhOJijigXiHW/k4fsDr3oJKgc+9GvwehsYYYEEascHC/CVJjrmmjMLB5kLOjZz
R+LTP4+rwTJ2Bun9eZaRTot4Lz88kTTWDKwLwAJr26EWetYqxS1fN3F/iInbtRHk
GdSVYNohdCE+bgrcZXebAMlMppSmvt1VHPIXanZmpcpcmKNvQea30uhqBLPhR1wv
m5XZk71Y0mSmlAXfH/lqEiGQoE/Vz9V39LL+9yX4UfdoZ0UXRFZXeJO1m5sAG587
pPhgSGSW6cC0sIf69725Ev2nh/NlqRWjEJmVEIcMVBHgeaYISlu1/YozoV0hiSrN
gAUlQim5itUQ7xGbzj/3vYAyUf5FCsmOw5IvCIc8uldhQwt/u5fLU8X76zyd5WF6
T/MxqMZbCB5TMBMLZDjy3pPdwbiMUF6vcIRtmtAQpd3ekabX80oK2Ydn3CSg+Yrf
Xd53HldSFmq+nmxrfvFFl/k3V43J1FWd5TEB2rzfZkRqo9Mb+GRhVSTmv/gl+U+m
JgwVqXiUsFXZrVqPBwG4Fgxi+Q2Twv7TAQb618VOV61gFKoQkByKbGbBLBZUEDGt
bEaK6vu20++YniMHe4Wpo51kfXmR+D+3s6GTWLdOnBSm+gVFjnp5+RN9e0MmiYjU
Kyb9QHovZ094yIIcJzsUa5/P2qDpti2YbUYhEQFgatQbMNCN/tofW8c5Yy/s+rOT
kUkYS2d6Ne/ng+PckaJvFFXKZf7NAsbuovXTevsrxzpjH2uvpfdXq/zvkgcjSPkX
MQ958VcjMAvqXLJQKxWrEIjy4qUAbMY+E2P8/kZGm0f0l6R1IHyz3E89cRZZ5niN
kJI+rNq1INDgDrdm3vE9MzszNpPs5aD/42sv2d3WI1alOlTG/tsf9q3I0enVG7uz
Zymvn5iD5StBIRTk5w1Fz9P5CuMf1RlcFsrohSNmu+FnCSaFKWPgEsbzXG6k2VUs
QKu+15LMPU2p1Pv+VqbRySyn7BOcz8tOj3OBLL4Ly/WmX2ewkt5IykXKmwfRTb3m
nV1Kv57t+T5BAlreJH9AAJv7BTKTIJn+d0CI8uwillOMBY0BuQ0h3y+NTRSz4fmR
IN3gWaMIEPMZnCFwv2CrWJQUsJMQT+Cr6YCB2AWxAn8DXrLXQciCc23gpA03LHOA
MhcI4UFBd+mYcRc8QvBpWnpI+6tFdir6DOcgvJKRfYs=
`pragma protect end_protected
