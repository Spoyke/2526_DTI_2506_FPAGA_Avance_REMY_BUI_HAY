// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZBZTou0gMPUeNsnMZlvZF5eJTfyT13hZhfIcNYfmQJZ/0+V+ANIKH2KpUf05Xg2hiH7AyATjok60
IP+OJngs439fU6zC8HK4215H+8AIlHVC9dKhE5M8K2fuR0Di2iZR5bH8lwcYF9wrOSgm/61B87v0
BYwbecE6HqVPf3XH7n7D3zUiq8sYP1HmvOHVuTEUr4woYaNPUAl/V1jTS2M5W5+WB4Goyti09EmJ
XbZx3jW1OZC0U1vmctwSbvoeh5cenUms/OH9gCFjoT0iODN2LZu/9CxptInjQ6baIbxyUl8jNPGh
jp5yozfBa73/8Ule1zdiGvnXbNWM7foQ8S62Nw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6704)
FRio0ppzqezIUeX+V8F+bHdJukLRng05I7MU4yXfGNJMgP6GH5XGhHm8uoaW7r0Co947kbyxGF4E
kGhsneQ4sU454vxp4cmExoLu+hOowjDFHvBsCc+UkH5TuFkXo/eWnjpz/RpD4jARcIko3YXFXTQs
ckU+/Yp3zB5EYaGJdNCZ193krytan0V2qxByySTffSmdRf7I0TzHwEIb/TuQxW7j0JP0Zb7FC72H
Er2bIfMtFNA4CUrbo1mmI8I0Bf/fcOw4QNFtPHgiQcycMbdBcN7fEDuhylm2jEul2UMBqJbSWz7V
bEWgEV2aa7FljRu7xCQ9WhH+yuD2RWi8Ie9i0mit36TCMXHFBTcTMg9Y+Q2YsxbvWWNShvscdJHh
T5lnY+SVGuA6XXAyFN5Dgq9Bwc71it8m78mX+Rzj48ebRz0sGIgxmeTjyp+qYv31nHF6pXBQxsLP
bqkgudExpqoCWkUTm4bLPKsI+irT+jLSAk3R0ZryDA86pVPi2ymC5X27hp4bM2Yr2ePRHxjnLDTJ
fMqrasomAnFAxe7F6BgEduPCtte9Phiob+ZZgEzMPBy2pTlW//TGJkTdgOW6vU1ujh+ty0UqBqb/
lxiXFsRMMHrZ88d3aua7TeNx4Um/afF86xm6gXAA2LbJmZ3eBEBfz4SuX66qRQOx5vC0VfocPDPU
EcGes3+ZOCudvvOSnvLZoiEL1F8na2NFmd7gguoxje/EYdc1DArUW59XrezL170tIUAiKj3FPFwo
05H3Xnhl6m2bGFzXT0c4+5FB+cnKX6iIZBFnAbMdvsuPX3ZzzB5bj0yqLwbcWemoNbVZPA87eEzl
f4jxm9Ga+Mwam5/+qrGB8CLVw/H/MsE8IHJNSDzcGk4zw71O6KL3XB3DmPHC4lRJT4ezyDO74RMq
oX/zKN8N3bNsxjZjKEVZaL7bqEeb4l4ajDh6y6NeAU/XxSmBrjiGy4++AJd2aNfN1dDNm0kNnEK0
+yRk3i141SfTaAo3o+EtsqUglpnI4ZSqOdN2L3plh9aLmtp696lpDNW+1/cPoHJeQ4BP7sQnOQDF
HAGpsKdy1E5hjgS43JejCPorU3EIYTsLvqLOirBAo3Ua4tETg19psIGYqOm0Rk/3cxarN4Ovts6j
6i0NiGkQqxdOyLvNfu/I0Nu3fuZ9+866WgMyJQwYjKp2BYY8rdxIgZKUZMPZpfhdtgbOJBDdNbYv
sLZb5cm1OZdEXrHbvZwpIIyCprKnT99WNAoWBIXkhsQGfrPm+lsAMQ91UJynZGBs7qlx44VAQsLH
Mio1CRW5qPjB+uMwVYStq0qv7lLpXdlyiqXfA8pyqyO3JxwGQnQER88AJ4QxYzHlLLOx9x/lNM7m
25BaaoNAxyYgq0iFonSLcbz2HJPIloERFsjdTm0U/E5qM+3qcu+3NDtG/wzHyESJkL7bzyGL19tm
CiHMj8qtxXxRvcAUjc6KCiqhz9S8bbMWkVDncUCLSc0hEMMtm1NYS7hBTeueQpK66likClRfD71Y
rRvsbS6sZEVPMwfdfP8RhPoGABwyfw9sIN1LpxZFZkf4axYU5uf1c8IF1u1rSiIigVe+WK7B9MpF
Ys0FNDFGB0Zd5rwaMJhcjvYGRUHKHhUoTKyrmoBb0s561lBJIGhjcD4qdRwQCHSlB6Y0B6xypLcG
hEd4VA6HIP+LtBTcHjgwxk0nwlWQdf1Y+eEehlA2zui4MsucpR/jMVf7/CtzIbHSmJVGJAprinE+
3nq7hhsZ+pSvsarcUAqQdGgi3hH61C/6jQgSe+U43VhTS0RZvTchExwjDzwcujMn3EsOnZxMGZhW
T2I7EaSx2ST7sJME8RHIwKR8hFvl+Hn5s6sKn7oPg0s7/bQAdHwkY6D4X1f1v3h9GO7Q4KjeTS1i
38Y2nWyDf0PkroJz6XzVDLsIGOxmf9UugQXOo+6NV2SMMgUSqZwhrxcxCq8jHte7ITOMNMjKfPvu
aXrKfu3fqyMIfnTMebi89oZRGF3+P44fRCZVgjskNsGJnWLDBdF3QmasJvuOGR9qWTvJpDNiAfXu
3+UO0Dfx2QdBIEmTGuH+yPGyy1PsCgFR1tOz6NNsMNLKlz/7RmXx7pZrKCUVjQsNwsdmLsk1jvYa
nhm9fxxLyn0jejJE2JLUzCA454bYMJLPuNgmAz7Qdn/QHT1qi5EIIBv21IdSH8MlQgu7FfhaFwRD
q4fFWayR5vlecXzLhdBYqsbWN0yKB9DxjMl4MoZEtQDnQLRdOcct16TYVSdrRzb/NoFidPnJTXFx
xbxBwPF07UuNRxx5GpboYf0Ag8ehUOClXgPFme/YwqWxOCILpba3a4jfl5/Bhl4fR1CbugHuXRfB
zbqBcleetptvZKE74QvLKlDd2mF4CTHGbmQ/ZwFgNWGJFUoe415XlJop1kTnXlz1ZJ83iOWi8gMq
ajz0RAaE5ApqRUdlrd2zf9YRGhCm314WLjShlpJXIpgdKe5KKCQfUDls1oNBXTp6ztPovlEefu4w
nusKPjJ1LUpGYcZb/xCrAhNCzOR0OX4+NuCrZpPH9OgSjhyft28088VEUiuFpDdWysIR/zjt94do
bj6NdjqOJzbqia/Pfy4itfzqiUwBgcZg9PVZZy/nma6TaojSe+mrX6jAIj3xc9Vanl0zzzAbfiCe
kTDM/AMwNLcJB9+WzsfzeYy9fVSSXo/zT3zOWy9FW4CEAi+HdcYEaMWHt7BQ7emASqIpFeG6Lxl0
r3s7u9PHn3SiOJfiNUe6LGHaYHWwPdTzHdVy4SQWR+QOzWZ6/l0/B5xHVGauuhJ5/wbHUqJ7MDHI
QwfCqqn7sayYFRea0z8i9PlqGw4GVLzJO+MHBRuiVOna2LHJ2LvLEiomV1BANFGu7ypdH/ew82YB
8EeXz/dXqoELD8nb6aQ822/sqv6QSd/zLgSOlOKCuazQkIHgg0MqC6shdr34JcwFwNHPUohKW7mM
SPyi+mAo7fv/16lT/5oJuTkpP7T1fgTZ7UBQ+PLCQ624DkRNR086qUoBO1BiyPjLQPrYnyrTCOjt
fb5ILCbEtj/flg6anJWF7u5P5PkBRX2ladyxsvJbXTE66JMMSfK/+lvq0Fnm+SitrPEU0Oc+QIEd
cySRCtafP97+EJPWA7IsaOwQTSn5luRl3TNv0yWi7KT6vYWTiqRDXdirZyKFRKEosNsctu2QhDiM
ahn/wxgQpEO1/3zzvmTJhfO3tHSbwfnXJFc0C/VV1GsQZHQ939cQNTGCwbueM+UzbJxi42gilhcL
b6b09nRXB1T1Y66fJ1PNKAUzLj6n1I1kPWdz92O5APbF4m/FlLeRLbZx0+ebGeR+PNo3h8uwzaNm
/maKOfDMzXqvaLJ3xMEbPBouDDONwCL3KL8S2P6xiWJ6pu9Ll1/X2ltAYg7Xi20A7fLKkLrJFj0i
lhlix37Dr7sWxohiTEcahr/YY5LuOTZry0g8VtrOuKjBW/EUdmFr3N0VpI/OZF2mP6MEtvSwa6vr
8YSXKXF9uCYCODQtgP+v5Moo+EwViw4xMunKI27LLo16YmmqTbEiOUdaWc8hayH1JQbyVmkODxA8
muBkgQVgDEm4OibhR0bzeY1UNTHEhEvkm1HVEHW7In+texioPYrr6CB09N70lX19yCtpvbLpBQUJ
MijAowKP5Bpr+Om7qSyq8HS1DgpMlQa6wojtIXUC2cKoKWD+wybrfXtlnU1j3VX0IeUWh3mQP7jv
tmFTG1u60vgKy1sS3b+TR5ytsXjXA30jlsG9ZETVQ7dIqbWSIIvdIYRjAokRE8VbCO5HuYmySV8A
ktLoqssgEY/vGsFfEg6sQ/YK3fADWuiCOTzJdszaMOvnO1h1uf1wiClh8LwSPxFjFfiCYO04KCAd
94ny6gnNdWheEZs1pnE6sB+WBTh6F6HyyFXFUhH8jV4VJhbc0pugd4CTsBLxhordGpA43HIS0MPs
t3ttC936WZ3E2yxyr6uDPSgRNm7lhEap8F9AHcr0EhgjdgJqvQkyf3kkmMya8Dk40oZqFjVkPSvp
BN82MNTpLjoLjL4dr9frUBcPt4vr6TtPfawYJkenmsCERwlaYV56KJ+7fraplNUtcmf8jkND8Rkj
ZUZ96dQONDw8lOOBD2XPan/N4kloiyB+0SJFFSVu8cRrZbPuX316LoiEWUcW/gaATiuZqPIxLWbs
Rp1v9OdVbhEnDEnNiSg5kL8rAXw9yKu9YB5Sc7/9PcfbKZn5qw4wVFUHRULOa+TsbKxS1WrP+8Fw
OwZN3JSUsmiBD/WO62Ix7m5w0pQDpfZQJ0715bSi/yz6kZwIITHD0WMbGKhjzMklxVB/xVgY1YY1
qM/A0HPuWtxLMIcGNyydp43YhdhLbom1+fDVUPAXqgv/t5Cn3aBTDdVAhVLPu6MuONlU7ekOgylm
a11k9P6EevMKRI62cjZmHzyiN4KG/KCF7u3TAJZHkDdV9pURanm2CK3n49lSNs1sy8CpZ4x7IPmA
CibmMllEhRQhsTNSRnHvU6es1tBebica9kHYfYPYkCTj+TIVnIc653fn/F6Cgqg62gONNt2CQUlZ
bZEsHxtW2Qgh1H7JVC8Fy7LLYPlCOGgvMWJaDvPnh+jGv6Fw7wXr/ukulgme9sI/TNP+Wq5YDFJd
5CRIHjAWrZeAXGtYF6+U7x25Q3DJLnew+yeTfVHTgA3PUThYCmJVCXq+VEezRlC1IvJ3PtkCTv6j
f9DuiT9eRRW42AhTdjjxLYyI5iTtDfYH4Y1VZDJJ2r0g/YXbGJOjPWviXt/K9mfOiCM5F0VomrlK
kzoskNBw82kECQZgkDPuamJNPp2xuq3/skOXWUu2qqNccoi2jGgH5c3ylT+/8QHl6ZOs9QgFjJt4
vHy58r1gG81Q4gjh8rCfovRYEkWTYp2JjChOfrgIq1cPy8ZINjZTht9JIyhbU05aAXxztih2Cfzs
ifceUmlGuXdiFXhQNFZgAK5IZyo0RlJHBln9OxcB7ogJiDSw+RCUnOLL6RUT5mqzuMwkCxhOamTF
bIobXlJYfsNBnxvvuwF/fvJveR422yxST4Pg/6C66ZUeaVCICfJTORkGlGeUMrtuRmUrWvXUcDnH
XAfqtRkYuYilgQBycwbXaUELUFFc9mSAQS58XsdsXfj4GNTXaiiHD7Tv37t7AIamleg7ZmctAEvI
EMfjtd004SfPMg/PXZBriQ/gn/AqVuQAgBk10B7FbmU/KBi3Yv/GFx5fgj9CBIIvP4jVAkHtMKKq
wNl+s5ZTR9txG7jM2/ZQH0aCucgErrnRgj4MmEpp9YL14hEn6rE7Nz/2SKwde+t2y+PQavPUQNGQ
Ve1RSyNjHTvR2gmJb8/T2hf6elPWdNHlSO6y2hVm/JprKPraq0BF+W5qym47BboMoc3kxRi4hOMB
maAP0Uga1Z1wsj0nX1nxiy2dsh5mhq1mDCS53kgxOnjkkmSNaat07s+J7FAnEj5owDVY9MPaH/nF
5nNyNdj+cZ8IlCwlzHPitHpyiqWaxb8Ns89uRqJPW63Ia+1x+Yj1MTHtFnN4zWqTGUk+nQLIwcHi
jNoWtf8OKNahFZksEsIlW5Gn71sYAXYXsX0oE01DRwDuTYUKhdN3vSjF2x5AoBekv9HqX2y5befx
GsnUPF7wXtAiJYoersEsgDiWF9pb+ocpS8ct6w5u2p9v3s1UW78nYKfkJZl2Gd6M6okeFZQ0J6MX
HRtMamqGipRthywcDvFv5MBoUHbyIDsL2EDfyNabhgaBYXM8z3xh3VhymooTUc/AIwbs2YfmACo/
2LnWaBl8NmjXaEfcteuLm6D+IT19/LA7miuPOTYYDoWotM+oATqn55ZTwwWR2VkMmD4bLpjPBD/w
PIAns2S5nB0oQlX8cT48pNUB8KzcCBHFaOKQ+sQoT7OryaMuCFKETuQRa1S3y7WuSKMHg99YRmPO
0gLetuGf0Q53kIOPXI8YAZI3nwZ6bGWKXuPa0VLA4XnQhfiuV3MSeMiTov+mXjuqIpNBpgVFr1Mj
FWd+8oxLMV9jR1Lrh7L07M0JCK0EFqJV03YHDlJriXdX9nfLukM7dnH1uylqe1ddSBz4O6qWs0rf
YlTer9FtlNRTO7Tt/atjUb5NpcMHPa6wxQ3grwan6zzwACVciEhzB4AEI29HGRLfZjyxeaooCzx9
gDs16pS4qoA2a9QMogNaDnu0/0/1TzmlvcTjLJ0CiO1pxaLGMpEVjNCGEMomLI/eS1EtwYkkhKqL
OZWtwyQO0I9tUnaiaCdMnd40lpobIbaHMatpMLGCOxCTdCZOn+178xaE8VU7CIOLdypfSmgv8UbH
LnxQfSQt9TaaWhJ0JhdRGo3v/j5xgK6a7q5za+VSM0isTNvY6yQ5paPYhQDgMUpIPWf6pjTXYcyz
rZGJDgG1alX6L8N3zLRm/c/D77R6Rdd8G2QRG01bjt4eoYaUmDI+6Xk1WBvAudKpwrFebVrzhlUP
LvMNzrnPmK7hdE2y0elcWe3PzPcudyatYMyW4icfjIg/fz1qLw8ENSQ8sfAkeIF4nmATZggYlOBa
iNWjFQubARM4gcl6EUFLud9UNd94GFFSc/Nk17nVl8XxdIAqqNFPrdkho4JJ4wNEXwUblbwAPnx0
f1w54rPcBYkAgP7pp/laDA4lUWQsI4b1CTdFERfys3RhHosBVOQhyY5yf8YsCBbVmTOic4zNdpZr
mrBzM8k1p9t09gWQlLrtGQkosN+Dg99gR7LM5nbtHOSxw2T2JbIFov/QmanHsFwP5DZLAatnC6Ux
sh5E5ZrGL317ImsxYX6vwqBypelYZ8fSO0JagT/C6KIv/B8eiW/FFEmeUGhMiBO6cNTNcYKIawP1
Quc7Zfw1te1z+UX0d3RWr5ekWFyn2HhxN+8muPKvi7cY+VqrSyoGzDb+PxPrBhTOgxsJDKD59kIC
/KAxYR7PUZz4s+xeBqQcMgezt1mX7idOr5PcSCo+iAtHVFFjgJU8UoRYIol6RnWBZhJXYRh3VD4W
ncH8BYCXcBlQ6ATbevyKjlgN8072KFxH/KQsFFZzCMcUrX6SD5D7YNsW5DVQTA3pwqwEVbyVZjHo
ihn4pu/zgbGh0Gz2kCxZ2V5heHoJR+fpevtLlMEBenMk812REF4Rz6q2fl7SueW9Rlv3EvXlf7FM
nC0RkFcFQqSZnJz7GhESMSNpSLKUgYlojDtYK30OYH5gwBIg2TJ6xR1B7MO14oQCDiasU+zfSYiO
vvP+iVNYYCwoLkSLOr98VJxn1HczGjRZloePhlrjdmDZQu51WxKuaAkk0lWwaOa9zpcRpGR8US+2
83/cItHcJ9h9Qi0DyEsqKfTasGTc9+sjXQJprG7yftNT3b5Zs5BQIlKCVhjhpNcZhFmfH8CR1ndF
4sYAh026ROSXScxGQTPtkQkUxUZrLrlAj9cp9Fb5VtbthKfDVr8N0bXr9d8wvKzvautnzllXLS6d
mardgbY+4//jnbtioX25hAtCmtro1TMhjXgRlBt0A1k5edyk4ooHPoeYh7+3ejw4JC9VxAiu4aQE
lKcQ3i54tZSiwUU/p1iSH/CeZsQM8Z43EYqAde3mHHgEh7eNLZO3vN0YWI2etlFt/ef034HJk4R0
adtjdwFp4OuCUFLEd2qGme6ZxIRDeUIKbXBYAeoAbdNLUn+qo9C/0KDHqbEEd/ivCGiOMNBE8lN7
6LhHNe7jsfkaKnkeAimuNa5xGGTdB9qNQ7EeX8N1XABi4Dd5aQpnM8Z9fH7b74C1Ln8ovFoHyZoC
2GW5cMxbz3H0Gw5zOTb62e7FNxr6nczPQwTS8mzXqwgNglFpPr652sLtsh4g3nbWTe5vVufduAQv
7F6udgdIwAHZq373oDHLdlvx11/ZyQVPWItKIDm0k1rTrbbDfH3zkoNDZkKdCl1YeAKa4esl2zNG
f3H0FPJbrBwhmmixD+XLOfpC9QOc73lJX7DmMGxaqXsIqHrRJQhrz9+GxukqSIux1tV7xkhCszIS
hJTonHrSJmqhLLYIg6G7974WWcJmt06477mNcrOFhlFhMFQWkD5Up5zcmSWyvInDPGzTkwmCRs1r
xNW1gzwh8ZybC27bThv4DZ8w3z3RMWvswiFYlqtM2Wn5qnj/jy6PyYvBxXd2jZ/S0HAcF1r+rv7d
pFY6zQlQ9dBHv3GCBMQjh4caIe/t7mRhHQ2AOkLmRSCxMX3WokKxk1USG+apVyNC2A03O6yvN9UV
IL2VWGtYptBVGCNlc42yP9sEvlC5vsUtxWz2XiQ0m858bGZOj9KmhTdcIXQkWzzpWIxnBsV0Jrin
ooewG6iI1KBiBb7svWySApVYZyz7mK+Je5pLS3x8w0v92x9Xumi2MljLvO8n1cjwZyVXDHUXLccA
7DZEahriLuxpii31hUZSvAa3sLVnu+NkqgE1KssyZPGWB1xH1FHP5uLSg7yuQfCIKqSLfNoIn6UG
UFpTFcgQWhzNyR+E8iGeNv9OFXiAc6zC6y+62LQJVOkvOJEy9KOFJmN+kW7MbwuD4D9Jr1YR7IXw
zafsiuToDIUwvLFniFjsPkcDXNxH/U4wE746+92LlFWLJA1pPJJxrKWi65BgnbEfBJ9TGDsG16s6
QGT190pwc3TVSTEJ4IT4mtr8EZxDszwClVmtp6Z3JKAGbjKDLHBgVlZptdSgDgQh0txyQJDXOdhQ
80mTLtVrtXB3vGclR11/uXvU/OkXaRg0NO47hb/7PNaloblJ93c6mHvzYtIQTfgxBln2tGPqSY2R
XtyKkXPWIgr9YADzrJbFVoHiJ6hxeevxV6sOEprG+KoednEbC7lOYm6XNqCezgWGK/4SisxGTyTL
FuLetGXFZtABkRyEDRxBKd+USfsppHy6U/RciM1mVvQ+2jMUPKO22n7U7Ox/cxYGlHLeIlEd6fqP
JBvo4rhHdG02CGrrlWOFGpeO35iFA2vaep3ka2PX1yWkMjY=
`pragma protect end_protected
