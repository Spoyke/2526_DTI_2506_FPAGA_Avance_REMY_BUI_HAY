// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
D46P7P9yMh1/3G5cvhwCHeXxpD1SHsNHKjuu9pbd5MyJ3PwuVGthhRx4eMiY8Wo7Ior/nOC0G+V0
HJDrbKU7khzB9ltMM8nbVf5guEW+k8zjpGmAXwCInsLixSYhLqNnoB88mkOM+JWeB5SZDIimbbLb
VMB2Z6p7RWIKRWgZuVW3kd6ru3rZH98QbvNg8Ni6D1lHA73NawMg5shLtAxwq4gabq65LPHIGgKx
+9GPoXyUacIgNG6A6ZMQYYY24an69hFEsVZ3s6rCH+ItwuK3yg1HU952Y4O327QCCFAkEff2Bxq/
/0hnomkbp8bBgAB9uisN+LvHQn7WQeLIJzE7JA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8816)
ZZgs5n2T5Wk508VGmp7cMvJI+PfZVvuiXRoqaDE6OdmG4n7bcPOCjDZmYTIzSFzlbcZbrt4Q8ySr
9hizbKtgzLUvzA1UhCuoOVoNiXquzo1M7J0o5BoV+PSJ0vFV+pfwKVH0XliEGNi95VruGzbdvHXY
rw5VDxBdgWCGN7ZBZdY2qxf865IYZtI8YUWmjiZx2NDCVEmMAWnUrMU5mdaFclbSZDl6dFms+Fyx
cOwZNeD5Abc6FSwF9zz80Rp00Q1wekpanAfXLnLlYta0wIY0wwDzhq6ejdF58dxBlceVL4nFrp3I
/RQqbzOAoEoFB4dJlJGfvbWzj0DuBR3eh+1x8CWKjNNB1b2QG38wxnBl91CXYmaPLhyeNzyH+V3V
iz5fuL1Ij2k0lwzbVu2gp6Q5S3RPaMOQPsL4iVWf5aWD/5VZ2xBWso1r5lu0o1qbsU+647KgX6a3
lCf+cGzCJ9mGnnfGBbg7Ed9DkVsXxGsxHGZbJsryPDJVHAJD/pjTg8sToMAQvA7nfgAYmYNZ4ABL
VI5GYDAPv8+HbqzEk7T7amUTvui4nRZEpt0niiBig52+6nhmRnGB78sbipqDXOcOe3y8LhT6xLbT
i9w41dlNes0AUFiwCjQLeDae2LlvDDsKRU+KNSrw3J69mhu6N6R5iME62IdI4Hk9c5MHO+DTyble
WwE7eCOmXYJZYzWndKdsyGExWMM3GYFtjoqLA/J9DM5gq0FTNibGLtSjafVO4uo9tzJQ/7QzN7pq
SjPNsFf3LfRYFWJ06sL6LwvzLJwv1PV7mqm6jUMAD0Q3yIMIe+hfbhO63ZV/EqLLkiP3ijVPSVp7
d0NTIEOA8R3XCUxMZSNmGheg4MykdYPoNCnw4dkDT40hudKNNuz822az/ZklqPBDGXtsPzQ0JfYu
KMc/xoIFfPT7Tjq8OeohXsE/dRVJ37VokpSG+R2o1aKIZGU+L3Oa7z0D26PsWrJSxpgWtoX5Gyr7
k2mjAv+1ufgmjKjfZbbj+nJrPpGrCOc0OyPTiBFcPtZDLVYMrqC40HyjEa5LT7X834CrIHYiG6U3
aPyzJpCjKPgUFMDW6R//Gr8Wixx+ru3p9MxZpr1FNjsf9mOKi0zzCE4nRtqG4fyTPCKpaXZhgvyh
tEGgZ2C+7AYqTxeM4jc/J3VMvT1xf20331Y0p6E6bmYNNFkViDegGQWUbujrLIbOJRcu07ZbbP+9
Xylm+w2rzW+gNM2atEBpdRd7k89aDkLXJGxln63zOAMLS7siaDHUrZGSXrUncs9z0Scv4n67vqGk
6YDsDQPNeQmpUKTsZKXkgBeb+ig9Ob2TJmLrrbUbIuZZU9pE2odW5jFHbXL0E1CufIfuHQxzLDy7
rrXg2bjTQ+q5D1iBRfDxvXM24hRjNsvPKbqD6sIDYyd1RN94LqJgGktPLZs7LoX3x+kIUmGy/pO/
5PlHDPD3EP2Leeit0ZRcz39L3weK9YZ8XHAS/LLOkEC1dvGwd6cFnQF/KnL6gAWFLnCl4720E6YN
b09MNAugwmak4/GLBYLipdxEldE1PZmRdFdryM4cqbmuvHpnKGL/VlZWtgMbn+jZRIlB35RIccGY
N86bosKm7wkAsJ8ex+ww65L2686Byxw28U6fqZkFstCgJGYZSGcnmbAUlcGX63xbs7Hj3JopNKCy
GWqck33bYO/vGC44oVdB6ZXb2ppMvIxzGevdd0MPi6/0TSRC1JxGQlDjvXpCP0YmeVIrSobf/VGR
3BHQQfEnZTyqXswrWDp75oHCbl8SiOv9JCFJd4kAuC5+wBzsF1Wer7NDUiAJVWD3bDEDP86Aye0l
YRo2Rsk/16QlUeongWkkCYxg/HR2LFmCbaQoAhIwEHHHb42GJPRAA4KJUyPhSggXF8PgQ4NMf/yD
JaFEKiMA2o7OJN2kac3eKkskcpBEgxi/xjTM7U1E3dh5MIJEq3nZ0+86MHS+0IefwKh20u5VkHYF
D2sjsJyIo7fRpmkt3rBAFJh/NOyB9Lo4J+FhCHSA3EZ91I9ecK91yjIk/PG/9Ia/8gizD3XCiefr
u7bruM4LKeCEJiFXpSaO2Z2hT2igH3gAOfd/XaqKkavQvxLkclEWa0kQnxBCKjstAuG+sGQOvWHF
i+WIesnc9/aIGnlwZARtGLmFRuNZTdg5LrlBPi8/gIfAn1xBj3Cp4XqViL5WTX28X4AByvuhXy1R
dYpZPfz0rzm3tJ2BvEPG+MRr27fNUn+k8rBlkQ/0UVPi4nNLVErXLeOoJrEfCS7sQ9rPf3XNx8qA
SSvJDhwwffztEyMXoX1soGQpRXJwTekMXMQCkn3jHBxzQMNIgRtbEry4CFGFCQlPrhUZIFxy10+3
qi4ER88K8lBuMUjh7IFFV6kfB2FrYzdpENPG0WafsvmaQoI+4w+A+EzGWZWR6RmnJpvrlZbgkITk
Tbjj02uEfuatkzzXsYf8RnabqvsPImgFEwaQI0/MyixEDBocnFJF4j+/HmFCgGeRRk68qgL3+krp
5Ff7SWTtp/cXhM89ebHoVTvbY4Yr7wXMIxOADamUguT7kMHFvHGdDeu9fI+yncK9nuQnFU40+qHF
L/9zwLGZWHhzRKzTW4FiRG+SftGKsaxBUtOZA+NoJcdLDXXbyBRGWYSggLFr3aJ+DiAWM0UJ0qPi
X12q2sSl4kdtszhk/3av4YdQc7zOkcB+gPZusyDVsS45gcFC0yF8+ThliBpCRaBYNC71xjIiY3F4
0Wm6SH+Pk2riyEXs0iF8uqOHLt/1fvYH6Rnbdfm35sOhim0Vogye+zDKp+WeMEiT3JbqMrlBGkuo
4Uu56cQIoFEoaopIKhNIo0LsVWH0rTo4f2iwlcEFzKLl8K8RAHqSiZve4lybo9Trzqd57pG9jNlG
C7LuyUHyWiF140aaBDwi6T3ZCR46sGPwj0YFBkOolNARzXkdFO52g2xvN39cNK/tqRKWTQyEwWsn
+l6iL8+VwG3co9J8jFbJ1cnzsr2bOZO1FyFdBnr8z6Bxo/lkdM8PKfwRwA6NjLaBZJBemhG9swr5
dsLszqLTf9Bqvgh2qRvGgQqSrbo+9sH6T/8vfbIkgOPgh1HOcWXmfLIaUxUCT0qgaAiDObSLIwPP
w1OsridHK030f0kdpZPzP8TheZbFNxMR6VH0ZhbWnF2Uf4BCLwEsSmzXCMcDhoHSyM7bPdZYiJvk
+RijNUEMldmXQ/dM2/HKDNNSGHTF1U7RWHmGOCmPMRHIwbIad/jzozSN3vQKhF+xl7rahpp3rp8z
kP7FzS9HurIsYTfnafWRUvsaN0thrgGOzbnN1SP8/cjV1IZZB7IAUxxSlh2ixC1HlkDLInEVeDIN
0NjRV4+XgWRgqX6AGCUfyy1oD9LJ89y/ju3+WK35kBdK4aDLrQEW0scsvE5A0TvJBa5EFlHCc2Cg
nIGpto4uQ+NJwQ3jx8wD7syJkNlehi7aFflZwuY4z3RwtdVmcu9s9GcoBN4L0ciGQj8+4mUowjtM
4za/u9H33Zs5bwrptHf+18tZeKMTcbVe75w3hFK9ksiIDuwVcdPjZeYWqJXxke2r9e5VxO68pzmT
NYpV1pgupTOC6tPsHpaOBa7EVJd1qjq6Ku6uA5tacadsbSPahNAm7r5B078jFMrFAhSU8f7oUuTE
dw2+2p+Y8flmjdFpgEQOuWTE/GIeD8fhbioawVAkTNzvzxCzQzjEUAo2hcXhWduIdbYMTfVtXhs/
zgFR/32LdF4Zt+ytRBqLfM6Tnb6Q2LgOvmbWqsMjihGqSU760LHYJQWK+OKjo/6kwknnDpfgXHau
a43pQ5yRKGRvG0C4ubHcTbN3yoWnMn+oODOOUNDRGH/Pf4nGQ0pnNXbhLDQhF6CGCh6vPwRpwk4r
+fAmTwU4N36wndF5xqFvIoLz75nIWMU1HFL3bV7hT+XFrN1j3sB7fyzZTR1nPeaRzghpQmhBm2b/
6m1P4E+iHE2J4OoTwR+688n78myfxB2aHW1XJxjExmPFtpuh+bY2dEGfr25Hy9ebwTGlQqMANAts
wE3okkIUYCyPNDRfGqWR8LILqFhtc6CAybXwVltHe8vxgbkebZnffwr7dsEtTREPnOtQjqdEgGZU
l2MOut9OdMcX4zQXUq4qMzvfK8QPBX302tDSdLyBcxzX69YTgKeaDBaLmRwvLFM8MaobRzc5YVWk
Qkipi1rnHtXVglxUhuCcGufiL0OD7ZNwUotc1GxdzNn5iHonzOW3f0VTn0uBggAMkNdN9xw8Mbv6
ByjHpVdAEWocxW2mt1dfFG/KzWJetgv4abGCX8zQEArVWS0+DoxWO1KQaI70q0A6pVNgqC5BgYn8
SuJ+GYtiKVvNsiVM/WGRIcmv4gd2UwRwUEdhmgukjGtu3/6L40m3RlFO5F74tu48BLklGy5AgSDY
s553zMkpNB6HQu3Xi/Ykc99g41HuuZPRmp21P7GauPH5S61jgP0wZwuKidPd7KgA48oQ8OoIUTWl
G5lCT6Glk6/hvmevxTGCUYni+qOtIH8/69HukKRbvRC2DKe7WG1HRRfBpTbYEU3e+/NwEBRAFoY4
2oixjUM9j5IilPPwLeO81TL3ktyzywkiKFw7XfEdtsIKxzvntrnANlTh/sGo2Yugg1GypAJGXBrR
jCQfv0hGU29AeyvQOHgygzZVQ+9+OEmzxUDb59dOKUnPP6zBkRi6J14kPLmOh7HbA2MqLIg6P/82
F/+7UDsTrwV8on5YRTuj731Rz0eemnL1IyfsqWssql89eujyZkrJ2SyWh2AQjXnhU1+djAqIgf9C
fewgfg5o1us65p8ppb7u8k2k2c6LLa929wDhOZL+To9XUgtSB5dv/ukfYYDCmdJve/OUKSqtyKQ+
NSyn5mmLrEqSVttEyQrIwEeEQdYAiirEbyKnvBnHbDTNpQzR+3BcjJsAxCgJ9fB2q3hDBwQFBBsZ
anKF7If2/YrCWbKGHuc9yjpo3yW35ca2uQeRdbNY47W+Yjpqlm0vNF8OFm8iuBYkXWefm1ULpCQt
spyI+7kkXsEHVEYpOMxTkw3DP5cy5nC7XsIfuyFMYPqjKFVsJKJUMAyviVvSSOXkePtgloy3TOZL
eG9aF0WA38vWXndvhz7wVQlQkejsduhv4bCF86T3OPm1yZzHCqgzVz/g2jDlqpt7zxXNO4uo9AoD
rPuja5+5JNZnxSYdrGaDA6U5JL/wRvo157CQsmZNvKLYt1xmd37nC/Ag3KTmatNk3bpiDDV4tSND
Vum6l+FzdmJ2haOT2VOCJ7HLtuHFHSBQud2Cm22wR0eIPf1BKqGLx+Icuzuiwa4e9Rz7k4alRmzU
NKpPAl1QXvE9QTXmDGfg2fEVAj4Ruy5Jp+U0uZogIUg5wn6NAAJAm5rA3evIS6VYR1zOIj7Ec4CB
dDbOvNMJc8FdH6ThOsgu4T6/zeb404UW4HzH/iRqeEKDy36I7txsJR+edPwxAL0HDoyES8hY8FlU
9VUMsRwqWHGc+P8vcw4Mw8Mcl2bmBpXatt5g+1MRXq/SQfayyHwd6d3cF3PUIOgj5wg4+vIHdyBR
RlYxvCw2tVTbBxMM/FIs4yRZzYPEskuJUURQBLVstDuwEugeK6EewjYDbvENOe8prv4/upEZ66jv
0m5n4kVP/HgeVPQj3vTRrv178476kK1RCPRgI13Qt995fLGN38pqckBnuVWUTH43HU5qjoNmssVl
ew3q7N0zrRURAmAx6nuEa67iSrCUcfUKHKm0pjItNjXw/9qnYkVBILzIeXce1nupclL0/7pmVdJ5
IlA2QDuG43hQQdhZA1yAUpBrwqNVYRJ69HKqlVKzeHLGuqkHG4vJ0GfiHWJRDqv0IkjfYuBaLTqc
emDNmtj5vcOoneL2xjQFaJDseaREKZcw0TDLTscrPFHynpRYBdJiAWy1648dditP6cau52VkBeiP
61FFfkTp4Z9mZxpvuCWMTBxxWABGZEQkd2lw3XWEa+GrwqeDOmpo64WYUwIO0cOGuPjBuy9rcT5f
5jBk2iN50tUaQehrRGxcCnYOIktujUQoefxu+PCWh59KOn1evYJFnwNC9mHqf1IJgWgDvIVbqLNN
r3xoOCDSDwEwdoSrhfN2S3Vk53w/eaHKDEhyz6QRapDuq2LYEy0LtSfmKzaiFjJYXDb0xRkIuC8R
mfF2JT/wdw6AE+aJf81g1klTcUKjrEj9XoylqcZYOnzLY2cxMWqABF72Q//QvvvYWdc9kJt7jyb3
ZVJCDFp4hgFfSygGFXv2AsQVWdyJ3t4e/XS9UYeuNEtVODUk5d7/6jWyQ8IVGoXXmT4Y7qe3bdna
0lHol6ZRVM1vyCQ1HpDb4iNX3SEIUhyYfIMymgjkGiiPiiYMgf6xNEgmFQ9gbKI40ds1yPFnrwSu
+FETD/Z9X8Nse8UIuKnw9K30jAZOmoTsyJEsDerqeyaY10krHMlPpI2wpTNN7/uF84JV5ylq1q0D
1+DyGTJukGHmGKqvJ6tFqznStH/nuktZZ4bKZxULfxdf1W3k0pF5DhRvbmdJKQccNkkkq1ZDyK5J
dwqWBq2yxtHhUvFep9OGvN6w5YkhSehEqB92V88Qo0oQpgIMx6IfC8dqZyNnBPYsVur0OSSzFa+Y
VGn6lG/5PEbIQ627v37KFL7raVdL//y4zEsxS3xqj0SBtkCv8OB8s/n9saaXoYgifnrW1Qtfh8EC
pGUN+4DqGeQyPnkBp+XYc2ylTn/UhTsPIy8l8P+ImCpsSemL5L6l+HW0Ib6qsYRfPNB8BmqOkKKs
2NF9z9nAoBBCIDPzkzi91O1IzkG99zxdWO3hjdCshWeJ+OBW1jC3bDWSFrfzhoeFt6c+0Or+c2z1
y1G/RQ5/awqQbVKGZbdct9aKoGPdrlYk084QoXHnsAzgWUhSP/3FGwdSi1Hf89FxJ7v7vPXu396m
t8N3Ox1CHfOFFBJEHH0Yap4++o3iWLbthPlMUG82YSxn7TUnAvoi7BZ0I5C+3oUQKNS9txJk30gN
MB9L7Kcup8+OuCFo8iqvDND5vQ8v5mYlpfMPsCJp6BawiJL/6qhrJhqW4XTP/CNlseTzs7sYzZ4k
+nPlAuLsUc2BVzi72OT73VshRj8PX0SnIxWRAGO0I0uGiviSRiA+/QiENbyrSDLPtxNRxaKSck1v
LhYv3Pxol3jwhPf8RemQb6VaYpW+JkUf+bNldZhQlbJLzRgqxw2Hr8m4qRCNhdJzoqDvy92zAKEt
M3cjgD2IMRJ5AZ0gBeJ4sh/c+q5r80FydLal8KkHS4VC4hCHJxCPlzPtrSsreQlydrz7r/S61hp8
aXXf+f+sHk6hrT6DYGn7DNW7/m/COYueVAgmd46bd8Z533fcJjS3o7Hf9ToyjjeQSq4PI8klE4i9
cR+k4vw0Qv3slMAMElNaH1ZMNp2iw0tpEKm7q+L+cuIRVOVK2UkhqrEgyDq36hyoWl/elrAS8hC2
BbpljXNJgcMFVB+g43/npQy6KASL+yl+S1bmSKhznXIFlMxhGf6cvbq4tGfoyYvUKSjLM2T0YUaz
HP97pE6Ak6BVOKYKbhH5WesNeCby2al5GuTCU0hCfZvqqS+KUbbSjFCyR0XrAUgrgQA44VKUq9t3
fyTllqsKfSKhPDiJVnfYIzZgvOIlIXW6/p6OG89h8XfiNKq2cNO3sgEcQLcA244O7lk81+Ub7cLT
ZhaBanixUdnAJ7AfAZoINTvDnbOdxAodjzMc5GQIzv93tu1f9Dow8ec5Is/R0XMhUfpvis4j0rjJ
LtaE2UWknQLiWVTnIXvn1JaK1r4FmzaU/7DdvNG8BCrhgIAarW+dmnmAUNePaeg9y7apteJt4T6N
k3qp/Lagm8SrzN2WwdpOPJYZc551EpQhCJw3doa8J+cLAWMDFf9CoAX1J7+lF9VANniIOhr4mVWs
aQcBgebAzVGUqu+Jvb5iCFCC9oDEqYeY4MR/blztbPgifeh3x2XY2OrAh1aNq5ziR3v6QSOeah/t
DOD4I/Y20PIl39KTsR08Bk4c6TTDqDT9PAIfnbpWvBBqGT0lBnViamfB7Fj2nctHOt09YMPqelVf
sUPrn9F7s7Vg4sunmn0hrrIgy/9ufWDBf6jo/cJ+x6xgUUiMM6owixkbFFV2XNP8VhihdqFPYFXz
IJy2eVbl2KngRH9rdM5oQMaqGa+2dhH+XII07p/YFlkYyZhI9aXDg2Bvph0NwNU6sqGZcR82Moc7
/W+e5kK4ORMX+Y/uMGNmY4uqaJkbGixS1I4mVjndbx5677dLwY4uB0ujrTmPXOnBqB+WrO8hWTKZ
I5tR0GherrFLIcLtYaiPQVRDXPIAOd9CXmsuwtWCF+zcFLBsWVc32rZ0gwsFMRuM9udFyoJRF7+X
JLSGp+KpHPfn/z/RALgQ2H5uJ+D7tcl/CALyOL37FIKYe6zPaYgVPrun0KZrYfTBCpdPC9DjOhox
a6l5awF3HwzCraYh55dB/NdbGsfwAFvlHJqP+STJ8Wva142TJvYwDU2d3Cur3E0Nl7oluodMx6UC
g2/YJGgC6lTjh2itMQ751Z7G8aLOSt61hY+Y9uFq9YLoP4PE53i60VEWW81kg8yYmexI2PoAToo7
c/Hl5gcKb2V8HFoMFHVUp168J2u/d2Li5wBDMqWIkuLbegj2qTGaH6qQh9lk/S3YapKDAUsEWGqr
D2Aow2DqYJOJKvnsdPha6sT0nCnCuKPghV7vNSnVykLSCebz4LTMVFzJnfoOksvkmwfCluYabxid
/uxHrf0PyNu4D0AD5npwt7T9yeAdXLuBq391zfbJU2zn32q8hAbeMTL9wq3Q5VeFaKI8Mq6Ck+Og
yAWq8KYRKw9uENMn+hLOWBzgHjnQnPN6vac7brSThxp6jvtBK8LmsyJIqqEdR8vhAa/u0gscC/Qs
N4k3HDrRlhOIv1NzKk/qhrIj2PWTVWOxS9K0vj8HsbBZ3nM12n8ppO+KaEw+KPX5QvkI7KYhVI1c
FlAjKkK1Z6BGsUi+NGUSm7swS+eBe89tjabfw+Aw7dfoqcikhglsJqULhdY7LOVJ/OAh+j7ys73E
in8tcuxEWlp8jdcqgbrxXIGFHeWxiY4x7CoFOXgxHk54XVpKE0gSE8TQCKRDVcmHIGa0hcqLFGAA
87Yq3nYTcIBnsDMTanh341uuayXajV4EkUGZzA8rXrIudYJQ9uEuBE6TN6rGMvOL/SrDMeqS2Ehg
RGgdDyrXGoLMM7V2AW+Wlz/Ci9ZCjoWf/sLZvFk+X1vVwpPyHohrK0Rs46/zbJuYuxamBuAI1Yxh
JaG9UG6xmEqHXlaQCN/tHFdwygm3qc9v5YCKn7MgZnsi3qWrJRPRZhTXM0Jgyi3JUMC2Jm7wwFTV
Nczm4ohaUDSyQ+a73wZb9rGjX/pBgnmSQ/cUTivA8xETs4vtdf+l5znHFkbbzgA3ViABlWz/pDLB
ifz/hPmU4+C5GIrxEERJR+lAkKvEAjW9J6C9qoSNvctgUvC56Nfyp7IgLtq1q+/YhiovpUqQ+LUF
y3NwkroXjuGkcXZsNLz7BxGQ9FFYHhgK1AIyJS0Uu2o4U0yUrmYq64OQ4+xaDNa9pAtYy8nkneE9
P+jg6Vg79ujJ4mayykvkASw9d3YRuqOOBQF17Tsnmf3eMzk878eWcSSYIchRMnpeU1KGjiqoCf2H
ttFXVRhzDuJpfii06/yeLAjd53ye1/SIUyWXKTYsyHuMfiEC01EUkXZXmzrQ4e3OTv4KkfxcZqB3
HsH6rFS+u1JHNGdFKUXYArri14WL+Xki0XuGr2zgyJsfneltxaZ8YqX4p40xczN933hpJoxdSRB1
1LfBI1c0xlTZU/drnc0D1f9STISrhVPIxGzfPVxjjizN/QMXWedfsObq6zB9uq9Wg74lO1iv4m+p
WUMLYlxOHB/zZEPcHJuXTi1h6EE+b7Me0jCupb5Lo763t55xKiBCXLmvsQHawg7Ik+wm+2hquweb
RNaLup/o2+wjYleaSrZRU33rdEm7jNiNHYJjcszKYVaPYrBSeneu4wnxZP5ho1S1Z3I+lT/oGzXY
D3DsI6RcPWgGWX2EOkCIiT0WEwH1wo5uIY7Z/fWt+OjZoi+zj6wM5SfhfIMKUIIxAe9TKzczjkJ2
Ah7mAAprDXni0s8Ly2+/uBlXYdEXZu3H/QTWK/is68Doh75aJpavN/LtsGh6nGDRUOK+n84x+KKE
7rVFzKrhnddNH078iVdMRYd6kxl0tERIwxpNOFuce83V2O13fegoiuMS0/AB6/t9Xfm7LC+nhGCo
o9yVm+8umxPmpzwYibftBNnBFIjDGvGeun3MYL2J/ayRNNAlEpUgjCivCEwpHa8MDDrWsjNvJJFz
V40W51gLBVkULDd17TEuKVwiK5t5wjRuSWyWkvb64sCRcoSwHFu+GANkxAuRT+fiUZYvXLYBzIm9
FfkTEndpjtGz4MKKMf6GyTtEmQ2byia6upJgnJjk1zU6bbbZXtP8GNrAPSH3Dy6ioR76nbu+dSa4
QdtHM2ehUDxVzclouDA9orZSnx9bOVx1ns3P24+zt8GU7hqUzjPaoVRI09NSM2pVfIof9j2YWQ6/
6bMTNfGlWpeFnZzTS7fBPwwCJmTfmCrIafG2KVTMoZpD2akQ5BfU6jbngQLQO88ycYgn8pPm9MvM
PClI8GzCzqzN+V0oWZ8z/u3NKWX7rKG7lu5i+H7XvWLYItZNM8cOufoA/YzvLUEDDjv3W2gZwqXD
Ph82lCacfr7zAdqOmrj0CJLnbx8wNGyw7vZ65JrqsbJUbME2fUQd9bqi6Dix5vuMjMdQcTPcI01E
AnMWGRwd0We7NK7kPYjSV2SQkMEr3bqAgkm+20kCGmWyD6Q9kDJmdQeEv0TbzJB+nEXUwDpHlxKI
/+RIV8xbt7gLY540zXW0HaLHcvaJ4AD+JaRgiZr0WeTiFHML4iA/lSONwErjLUWZ2I5aD8MR6x1R
daAumEOV0+m5PA2bREUun8MI79RdojBjc03czT/NpRtvXzLh0t71TLtwXSXAtA0UnDsO9rjnDCUa
uLYwhTvQbqxLvO8+viXOsm9uD09F4HdQUXRYePx6qz3khcz2jjPmMrXXOrcfaCY8aJTDNRLJK7ZU
JlZTUDR6FAp/UlgGswJJnOeLWjpn+QfsFB5OmIxLXy3+gbtRS8TgJTdG8SwlL3XEUaDcAgmlPJYP
g/Om79fpspFQxOzMhflpjAhbuMukGEA41jX7yEpGR07/06yqhg57Tt/fUL65VE5whbQQ4/X8uyt9
sz5i04AAqlvmlkkMW5aKYEDcX/4k81cEKHZi3vPfUa9v5nEV/75CiYMxDki8sEeRbAmtR5/c95N8
by73LzU8OMDJhvRIdYtTNWcXICmC1oYwF4HNugw2rPv0PZfMEHSwZDn/l1FAByT0BCLNYSmoDixx
/6Xuc5fZWVC3riYAdiUhdE65PuEHdwozcfDEEaZL041B/Rc7Kl4+vbdcF8V6owyVtHjA4bLozXvX
6GwWsGQw3uW+hngFpSukxUayOKSCnW7yErtGKXk8h9ZgUzF1u3CFaoN/ZMygxNP7w8vGQNuy/fAZ
5rrhkULr+O3xiBQ8Vmr4ZevMs75xuPHMdDlrRfFDD49Js06GvAPzqp1J7LN1x05H0twhX+DOYfAl
6Uox99uk0Nn/2Zh4ZokJRBYJ52wDA3vy/gVyfbgdB61/Dx5wfSdyjbJGW6CzGSOsuDCvrxa3011d
ycuHFUfdbRew2UVxm8CjB9G5ZnaiQM7ONCpD9rwfOR7vWW0KtNg=
`pragma protect end_protected
