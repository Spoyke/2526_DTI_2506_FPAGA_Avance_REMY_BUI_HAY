`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XPivq+Kr8p09Ogpe2Mzd3KzuDdgkR3BS+nA1xHk6H0GBPN+SwMbBI+HKKJAMBXjS
IftD4wlKoH2tpUB1xF+3QYhU+5XMlr/qLY63QxJRREAFHJNiMFhnmd882eha9E8Z
HdPhi86jEX4Q5yMfxNWN/o8zBjtZe8oqH6wkZWWKirI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5680)
KLpfv6kw1EbtRo2fPPemrf3vzGs7lDEG+FbNBBOrPZW9GC2aIo3QTCx41cU/5MnC
6IFNpHzRwPUCPMP3bSS9KEXkT2ka15dzgmnebhcTE8flznPdxRQoMEFEWtzVLYKp
09xFZBZWuCORs2eL+Rb3qe8XBigUqC48QmZouC5oqV2cgLcvFd7EtFRE9hSISK/s
+NGCDgDjigcp9xLuKcUuiR1HaE3QqobDh2JOKxY2UUkGRnTS0Ik1x7sRYpMEAzuH
59s9GiJrMi9Hl8yG3iQk/wKxI11Am2xcMboKH6e8upQgsDZ0dLrDU03NRgyKhMGZ
CUuXAT14K03gOZUiKtbK/HmWaS9cifG/QQ0KnPemKLTSeT/OtfZYh8SgJGRtikme
hlgiSoke0T76nIzSCoiNmAlZ/Lfbh1GQOfi73qkvItXe7TXIhnErkC2EdH5ZnYhM
ubpJGiGNLJuS/roD3n5wt/MYhBRj4XlDkMZqc2upExBeHRZUqWfoxHJkh4D499+s
YjghUxW1EBysg9+3P26ATBVQzxHAgD1EC8GImQLsqVAxmb8K9Xn6cxXjesl/Lcfz
Fob43ymtkMkK1SRTyXRx5Q/Jev0pHwTQwpTUSh5Vzwh0JdikxmSgu/tLkKLsAIKw
wwd6rKZKL4p9R0XS1NS7HE0F4aVR7bL0HZoRN6st4gALq2Jpvtiu5uWoAdirO6Q1
iepfovd5FB3PSc1/wd+S7co+AQ74Opb2PSQQz67oMe7Dk36HAAjwrlc9qAncY1vB
0JIqzXx/nx15mb3/ZpMQveOTTZrHP/bvHXtS9qKdopCQ2AJ61T6f77h6YTYVIRDb
b866UL7qCpGkpsHEe+7GWx4vaFMWvQLNc3aO75lKbe2SMSu7jn7UfZI9JBvYKnKZ
SvZGyKQv5pXMJSctu/P0sTs07xrC4C05HQYoG1Sks/Xg1D82YRPd1nQb2UyahHs+
mw8jOlUlgZZlVNSAhkwsYLSdjtcVVg/nSPwZx69clP7Znv8g18o3wknBDJOMorYz
ASXJp4oRTH9KLemdCgBnuH3pooZCnnjn7LMH/3FoTHT776mdeIYBhkWFYBdcr6pd
+eYWzHTmelus9iBSGHfbqIsh5TX7eFej9xJGlgQSG7bCRX+A9t69BR5byqCvxX1t
Fz+qFpQFbOIjJb0T3BZrKuavrjlC30Of40pxePRl3ZdjppM8wOErqzPh2N9Y0eWN
cjG/bHyNip4YbY0kxlCO3Lq+mb8uxUjMZv44JJn3iT7f6xVFM6MmsyLAT58e8lKL
TGPqh540SHptREYGAPCPt788wumEZMxVwb0Veq/EIEgjvxdHDLBUNEx5gF6spSfk
LxWQBPiAaBOztElCBoXRE42xFZ0YFxticEmIbWBfeMOlSTm1czcOG9xjikJ9Fka2
rnVf4r0J4cT51yjJTYkgk9DioObXkXI96O8hxJk45SGp0d94mi96xRAWsJXZ9vgd
YBnMhnNiwUZXuLS3SQ+G26uO9mklpUxyRApvjWFdomeeZJyJlD1JyWUx5ddatePN
uiavsN1JENzzq2lDhJJ+yZEe02ZzDw4qUOiT43t/0dsdrTD9/vPk3Rcp91sROIIP
DTew8upCV7g12HymeJrfvIenI+0sAN8lCGNJilDmaJm0Esh0m5L8HllvNtccFAj5
qlUakQq9NXWtNesFDly7NTTWtM5fWppg3v38FMmC/vN/hqsd2CH4ElBtCmx6+MYK
xUpQZ0GYEQJR7pjrJa9MYhLNi9BjUmA5cQ7r/0Lh7x/PIrdBEoakMsCYB7mzHb8U
s7Rh6ie3onsFeksqvTJXDUR0tLg4Iw1M9qdghS/DS/mfo0oH8HTfYE1m7pWwRopG
03QI2yKjSe4QUOWgzwnXG8PtwId1qURKD67K/TLgN/YqNO+gECkuZxNPesACZyoQ
QMmi6tmGvD4u464aRMW+Um5jfWldMvR2kPBiCpcsojwNOx2bw2KR/5ClHa+d/8vN
2KwrBDqGGkMijG10otKGxrcUsQK2LoJKqngr9fqLb8QujqzgzUw8eUsSemVStMZF
S/Jp3CY7n2E1ESQzHYRsh+Npz2tW4sUCqByG3BuRKgyXTh25Q/EgwiAlSxpBQctL
IqBo80FB0Xa/SFX8s5z7b9I0PCIS1Jl0bURUYQhtL6oA18ITqp9RiLBfjMfTsq+c
xaeP0VbUqq7n7I2ySnRaAO3h2S8a9Arg6sVkQVlPE38cL6F28eBjFiPaATvXz+Tm
6eEpdR3+rZ12sm/tVPTRZvvmPH9ULff5ZRGG9oI/Aj+Py1rGogJEyPZdGAp8aCN9
S+GaTAGY8kmYW/vXDh0XdYTZchVGl5JrEVaOMW8CyomNvpIx4rKEHg57LMOWq1Hw
PnGBy00eNCcztZwB/ems2AQXS1cBO8sLRJR6ZyBtIV8ChdSU0ucqTCTk92qTKq54
KlZ99JwNy2j2XAJpAGWbpk4ZSM1UsSh7jJdP4oSjsialayO5kTpAhjahpUh1KkQn
6I5YIuvP7fgsIw2hbOFWahmWeRvUU2TJY7guIFhA0iOIUOp5cU84Cobt4RQiuiLH
ePlJfL5i70m64M4Xpp61f7uQjlR+GtQQxnRsPopcgppZKBExUj7FRivDSBlOBXDT
ssDS8ax/jDB/K3P3NnXcu4t+P6DGkxcnEz0qV4gGCQevwkSrr2xfrawiFenTSdqS
TiUW+1OQ3AKhmVvcGIMKDK6fuzBqfm18IyTKetHMNIcoD5yeUUcZB3nEY8UOwB9r
LKtESeCMeAIR9RhlQ+trkyd9tqcJ31/QvqpFsinwsXZO13o31EPdNgfu1REaQF8F
3lF7LLxBsrFz2r+ULu1XJsEFhSpVhfFz3caHAqnhMH1kViXbdylu104RfFHzsAIl
3eZN2jdpWQYQV5SenjYU8T8+62YsI/ZGEYglhdqK8Jn0q1MtYUEnrFnqgjJVYEat
ZkqF8hJ6Wyq985F/3bR06Q7YL1ZvtrRhB1J23J6UVVeSjJ7tWS1KglNALuwCMp3o
Xd229Xaq9iELKV4z4825HaappjPpUCK4Jb1BKvbd+l/mMnjLbTFKVgrq3pdGWQEr
eOoARCmzeWk51cW8xjzi1KQgr/RPoiLk4QQxxHebTuuRAHs4B7atgjsq4s0H5zCt
oDfE8Z9RnHv489/fu0mwP0XRUldhLsd7Se3VHwhvKkyA259vMRPmCQHwb9ulqfHV
FalmzVV6qQo3lweqGluzNsqDWxx53CGRQ27rJaQQX1yXy2tkycpZIoMQ4XWp1hfM
A71VXU5ee4L84lgtc77Di/x2y5mVBv+4g244c8M0X1thwneUjzMc00biTBrklJoN
CsjJqiqqoP333dEKNUDEa6D/rPYJXrOvLR87cLyfE8qWB07FMR7dKdMjlcZeqDO0
1UaXSZm8EHIRgHk+aSvTu0HZBxgwxtV4fhpztnG3cO81gAehMGQ79VE3lZ+4CEIy
tRhONyhL14Iyd+2V/Qe5A5AEvgVv66Ey3JUe62If55i0s+IgGrHtqVCv3Wi1kX9b
VdEfEH5G9eqE0NQmbCW5302nOn6WdJvR6d+dsG2regLhs9Qj5CHZ9aryVDXaoIsK
63LERS+56A1zD2nKn7ygJexVreZz+P4FBP7xFVhpQuAEVr28Ko5wMbdYLuygfnm5
Z9/SATJzf72kPPJu8f0dm8BoRTANN8q8/xhyoU6MRnOIkco1XWrT/m+FCseg73CH
z7TlNX9yP5yxzoIL5k+ncUxxX5gO4VoU6OmT+63t5l6AI09ZOevC82uekqeDmZpS
/Kn5JGWk2lXSUiaNXGo4a6cCtNP62IrO/4/14BwVClStaRV5p8BhcRCrK6eQyH/s
Cfi2dMJ9oTEd1R2n07tf4rJmcr/ASy8Q19K74rb6u/yZm2nIZ8C0+rFurabpAhzG
9V9Ygxc9krUH2O06isU5bqEgal2Rzi0p2Ijd0wT92uBXOpk99l0F1gfvGjRL0OAk
vK1xjhiqUA92PgLA+kZ2+D5He/3sUW97TzLkSXzq2lX/FNikiM3dcWQXdEtxfCqj
BpRDZOg8LgZD5m3Cal68/b+3aW8cBQ5ED7WrgYuzlBd/EXFsSJUL0ZTk1Pim/y7H
eZ9d+zFIzDgS/ZkXgTo8i6ubbS/3E22ZFtQWKUQngOIsdQzKf43ABAdHbiF1+Soj
TxUJQ90xlLyixk9HSpaQSRNKZ/QwFsKugd63SLfSzI6QM9GUkjjHA/Ma0qNXb3Hb
rjmoVePHm+EqZloeph9Jr0C2RnekDkcBakC//6zHHBP7RC4eRXTiCnn4M56LRGeV
EcNad0oRlI6DHs2rA5OagV9N6pxx3A0Cq+97/JeQqEmdTx5VYPB2g8X80jI3SND3
/NssJ8838kp11zdoEqket+WETsFglCzYNi4myShDz81gUNtFf9x5ltKWEwxGR+mn
ok7MyMoyzs022ZtPkeqXXttF82IuweiPNiTurTngqFl1w7LbLLwimWCajC+sMYKj
uejNapnCfmfKjejFlYWUaCNFnPSzJ3Jvn0dkbZDkq0ONxgpYVU2pqBTwwGaobK6h
o3p3iK1xzfjYTQl7uidUJMw8GEU43FOsP+akizCpzIizL7ZzI6k+C2OYvYIMx7I9
8QpJrEyyotksI6bbaRqeSoxmGcCk4DMp0wo+gjYa98aFtq86o8vdpfC6WXjX8NyF
H1YhZEWiQvMFsaW+QqHzWhmRnU4TgyRqaa3w7SsKpL0VyG3IWkPCYXZ11LBITNxJ
PxR397ayYi7YNDLIvTIO/ks0xx8LEWZO/ptf8rWxhjRh2p5DkAIvgH41IOkqvr03
9s1omK3e4NIiOrTFTLb0INto6AXykLN9dtUCH5f9jkzgiZbsI3Y9YLwAQ7KPPP4B
StissZN3hnsncBKk87LSSICXlOMvWZ1aAGJqpMDVzXogmqttKQodx/Mdzk7m4N3i
mGS0WVCGv6dYOVEncgv7UvdEdP5iDKIiq8+KiACILr76ktfHVgGwI0QuHDQgZhYJ
/f0AwrD3r3jxuqDKU8mt8d1IjR++c7G6o22INkId0II/8HNfg5vhK6xIuCBRK7w/
Hpbv0+NGjMmNitNZCqA/e0IGfl8DOObjpK2LGpwy65JT5nhGIQFThoeIPdTZnkIW
F6jOzkKQsF47Nb/9wqqlThq4ldh+yTOjCYBwDW5LAdoLxQX/LEt7AD0TnP8K2V96
NC3mHwOJtOvHCMYtESUcKMwbZ1r2MIbfsD9alpiTDBJWHunD9Ys9Qe4l+g8UCLjv
7aCedpyEASv+UFdaM/ZcgY1LqM6k/sMcL4dPjZIa+fupWWsGlzDmkAdAtcbfsqQy
YXzBq3EN9vXiauwGj2vk/QJaj7jNhRIe7EcBAK1NkQmCV5NeUJ30k2kRZ/uj3XDQ
sDINHTNW8fw5W1l066PvmKjjGTiU0Ilb/LlRkMQppOwX8mlO5bwTyfnf6YflL9IG
g4zgRtmbxovfuxbLcF0Kw6kqvNlxF4RQU+3P5+4FjEijydM2bu0kJEouRh0TgvEP
rvF4ytnCN8MQgfqGlWLH9tha7vZzcJCzfWLSr840iGwasoVrIdR8NSOTmEIQJPcV
6pRw07qaBIzbL7xUMEL0BF2raN4qUnlN9iTdQE5pld/q6s7/jZsriR9cRc2u8bq8
HOc1Y8rnc9ODyO3ZOnPQKcPypnXxjztXltJlPFRLYjBsBOgUjTTXN7+jbxm1+XJ/
2Fz4+EAoEgQt8Vg3ONNlAQetfK9Udp4qT0lH6bzsvDL3kEBV3f1tZrYdmmt6TooM
Z0I5qac6cXDwAoEMSSdzAjrodheEHbu6DU3KqXbfa69bT7uFebq4Qejcss5DVokx
BlfWvHXBhaQ62OzBawIQHQTq0JZ4uZwx8wKpbO3P3V2eUEsTxLY4qv7D6gjsKabm
FqRtahhAiplWh6UH5ETUWtkFiZnsssmTbasl1wVRpnb03vOEXIp9pexpqkxKvYfr
x4QhmvA8bQSgqoEFfQM88+OxCCv3Tsq5V9ievCcgkGvle3TXBtkMmyumKWvRbQou
4feSE/tjtw1A4d2T9UbzYLgjeyPiXcoNhZhBJyN+KL8zRcD6hLNmehZYPc9x1Bdb
nxwMPuHkLG/35lSOWrYcc+cpKEfox+eOuy8N7Vsi5VpHzKkAlLXGFPO81NgjEIwZ
6TxNKZhCQdUsneABUKKfcIByepIs3EGkqSKYw/qSw3lrXga2GYCYsByHllk3m4XN
JVLkHwuPCGyUdcDlWM/03PoHwgIJQM2bv73YVA0TjsBn4kInjceN8cGAzMqKRcZL
y/Gv94Dz+Gso/JUWVkXmkDM9vzMyEEpfoRtnJF2FrNHHO+P9jiHkmLH8pv+2FEuF
Ua3BQQruP4Fk0Lxhjbv33GJ6Iv+6wrZtLJR6qnosoChReyAXPyxFbaB+ZbAsMIKB
u1J8qIBI19xEEFV4e8d19nBYcRLRHHBitbU31YwFcuVje/uKmJ9TgxKpqNs7WIvW
DUHeqOJCOmrK7LI0W90g8Ii7lQqRPhtqSZ18EGlGsY/JRIG6A4dN1q6HrtYUIyAw
radh7PFF2eD19CJSYboxTcc88646nILfB71qO3rg79Hq9o4aMfdhAz4qKkuaf+6B
UydfS4zdprrZ9epOnSoYfL6yUW86fnX6G+gbc6pWqpHma1BrmXm9JuH5FJunxZdx
ANJfsBZ7fz1nRJjWQF7X6ZQug3sz5idZ42Ln9N9L/0LzTXeKi3Mgptz5rkx+HAMs
8PH1xB/xiHptpdCid2Zo+LWvplEE0CIhqjQzaxPJDnknOJRxFiUepHn6G0UU2JWN
ESx3oXVhjlLnQ8otjQSXLI/i6beX5s2GCZjJP1/dMJss9Qemt54rn/utHslUBu6A
hJqLugvyy4FORCbaC9MCp0OkZ6y1xVFE7TUQMjoS5q9Govf8i1VDN9GBVzLVsguA
95CatbdZAqQxq9wN0SCAqG0K6j+x3Lfs331mBetwuwNsMB3YV/yJDv+/iy/5cm0N
H1iGy6wCq39dU5w4PEHUuaRVI8I7sznvZQUAmN1yHhOr9Qj6x2ZelywRJxv1D/0H
1T/zmcE4xKTDl3xVswDtaogVvJ+57l46t4ZbFqrHd/01IjgfCakNPvbc/QONFVzW
k7cE/jQvrieChiwt24bSLtshEXP5+tIfSdtGhrbuC47WK8/GNCdGPQhvBwxCSodh
Edl1rhyrw0rAlLtaT5NXBcQiWgzSXeZFRvqOcbwUGB7xB+bEeFnhLPZg5LvagIzM
oXudC8p66Q2qv5ywmJ3JQh7vKNIGnHBcoBvvREsw2azprqUO9qvKaNRBK8IFGwXM
VQ+g3GCq1GW/o7GNr7+hEPHPwkWoyTpBjgqwoFS5TR7TAzb09ccgN5JxfldfIIUW
POrHQhuPHazeSy9veAzd/LX/oUbYLcc8zyQyMY+sACQmvkCRTveTp26oIleTfvqa
TTHie2o0K28CBjj6yNk8Q42cDkMr9DECCegvEfbWZiajX1f34fmT3o0K4hcwOYjq
SKvilQPGaykK1u3TDOywdxyU/xa7+cAEJGYoGUqVGMQbQ/ORNG/MQCtVVDoDyoef
WAEuTAOEuDHSjMe/DLoBvw==
`pragma protect end_protected
