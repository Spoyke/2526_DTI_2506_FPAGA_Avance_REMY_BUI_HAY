`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L7BmSaaFXoEFCQecNMmR8E7PQkwa0ovdukP/PdoFz27+LLEdAejlD59TQ3DqlOM5
fHAlrov4uALX0nQQ1szd+ENl3pNbSGlGLInMMf0x+7lhYX1nqJedmqJw3Kc3wdmi
2Pu+nGE07d2zBe4xMkaDJijD70O97GAjCpepKQ/Q/Zs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7296)
lw5bwuerQe5EmytHEE80ORWtaqcBpl0m4vc9blB5Jb9NNi/u/oLm3T4X9QRlWO3R
Wv42WFfwfkA9FZqHx9WxXJjTmEyrBjPlHFz71mRfoBx5s2s4V6FBpTsJvWeauhDg
YO5HGv3J6YMzrxoYXNtsMsGA57QYAX/uojsxN/NjclDVIsd7Ox4IzzbgSMuIVoRO
qKNY4vFvdCgJgqcBiD9E3u6YhEgKUiiICic+SIv3TwkgC2YbSI0GRv9Yv4I+DlpR
Iam+EZe0ARk4lMad8JQ9vlzLSpnJP+B0gMW2F6Tsw2GCUH2i6Slej4ZJUaqn5mt9
+Orp1Sp1RkotRHvcUKbUUl9Z7juilFckojuO62Q9dm2rEg1lvkPanEhyN9Tgkhkt
OYP1m3cOQ7xt1pFY1eoVYA5NB+qnarFE5DpGv8ezFY1ULxfUh/wkbJmU3S/O36im
hW9hv1TiBLbXkJMt/Wpgv8u4WKzHGM8CY/AOal8T6e4v739T89G//YW2UH7Jokqz
vMylqg1dpxemZqSY5+66i8UOOAmn8ntE0dL0ntlUGGx7PDFN9ecNdqhaoQ7IuvLG
QVdt4YKzGhE/pfLZleYAQmZfLEZswPeBkpWbYwHUWiirpd39S98kizNy+60c+Aql
iDZD2SSjkYMJ9N9WCQlOVqoXZMHQwaYcUjaPngkHZ9824Ym9CWzn7PLeimRFIIqL
aa2/9oT9a4Q3dRHnJr0gG22Zb0YnsLxA5g1PgL2Zj0ZwDWMJC9ewQj2wyZXhqABY
Iqjj0LH1OKrrtlgaWxFsUNLH30+PVfQHpu8U+JTzZL8BH7+gQDhjYcUwP06Mcesu
RlWj5hcVp7ueVxR7ha10W6JskOm8KInUdtmlT9HqnMjyG81eYXprq/ai/X0xASiL
TpYseg8HF4YV5z3Z7NMyCMpgTjbYyYKfqYn5gNnCnvzhMsMGP6GsBPWubKXEN5WD
A6/TqgkH3hPJ20yvzE45RHXDg2Y5o+rcsqu0L4a0zj5yRAXpcI4VBI4gb9ug/NJ1
qxL75XA6/zHIFLJA8LvXOAdxXGipmpLx/b/8NmaTk1xqUpqwrCoX/Qzv60fS3XU3
B+JvtzA1OxhfKj8ohKSuWuifyicxhuABR33U1vvdz/pw+iUlIucq+tilIvKgDWC6
56PIZnO4aw2LLwC5AtqdioMrgZgUpqzxV0gFJEzPJutqiFl7G7ujGZqharrCBw40
IBFmZYE5Se5/X7jN8x8DrCwExBwyd/GbF/2vYS74pBSZer39xKWMGYQOF5M+xGoM
FbRv3sppoIF51OmS205ejh6Icp3oWi7xOY6YB+5oKKW1PmnIH3lhcvTYbyL0XKwj
ByHDzAPGxfG29Lj0PdC8Hbbb5wpKq7FyPDQH1FBARwQipxeDxorFtVhgdsb0PnHc
0LoohJUDXnBXke87mZSVZ1huw2zHk4VyETW0cTVwchYrVZF8N1yi6OZGMu2c41EA
b6cvUVev66nchvmr+rYr0BVBX2lGSGycVyL7GfX0MhooBff0GjNEH5H+tm2rhZ7q
N/pN5GrsGbh/1LjNPQS/ZrWl8S6sNVDVcvvzaZgVKr/VEzRzTqNf/r2MB7LRfHGJ
gKKMTOP8kilvhel71ysYqqlTDl3Hicy7sxP64xevr+83GdQIPshCjb9wVDjJHfLA
NStylvyRgO2U5+r48gxAMA3qaGcuExPChhpz+3GhXuFL4/oVN7kq2HPS3auYPnv4
VehqJUuCF4D4PoDfu6mvgk5Bpy11ZIZBkFJ6WsMpE93hVHAXJIxDEd8rLXrgKN16
zZ1kLWw8unrfJn+61NQKMvwXWdKXNI3nthc9CdbuGYvjQqkawjzWPUBaEr2ye5qE
q2KUpdq2O5mT9rgwa+qq4kOliNzOCW/yIQCv2ZyEMjm7yMAOHh149wJg4/YUT6j8
a4Dksj/lv7e1Cc/x/j7M3HLXE9LhcZu6Mpj9+cluulCd3I49KZ7PF8T1hflK7bPw
pO6s5oHxYqFyoK/6TZ1gspZYbQOozA8zZ1XwhaqQaq75/Ugt6yrj64ow6ptgoqVT
z3b/TZP0t+W7m/e9tlugh51SjslzONYIwVlwbgu7HcP+6pjK4W5tZcYMIheEKvi/
oEcjVXU3E+frXEdNUG6AD5c2xdftD/it6Sm2LMfdXvY6XBqYnguDXKrMIq83klqo
mNn976kp6Agcfg4DjiLPRkk8x6Wz+JkaMhiaK/b3DrM0fVZkMjE+tHHRkeCeAy8Q
xS1cGLbLMP9c/rijT2rsEo4kvIGQPm85UTBI+r6cUQFD9VWQD72IJ9P/ZSUF1DjM
LXTGoWr0va40NaRyYykmm1AuWhp4O2e/6lpu8Gr6z1TXDpiZRYp0+w/Y4EbkGNe+
wstGRw5fYJKmn8mlaM4BCjKu50ZRTGlErdz04K+7dAUsq8WN6iNenw0g28I6Cmzs
ed+BRiSYTZPiJJlopTNxoaV0q6JYVAOdGz260G6/nJaTTgbVjI2daqmimiCeGdLP
8ZybQbJVvTALkY8vYAq9DIJYF5Xhh5Wkjo3cnHdTI4j1er7SzTFrlpCVK2eNXUFW
ww5eFjby9A8G7gH72wluDx2AaW7EdatqGxwUjugp459SYzJqpfam2V68gKH2WgDb
47mInr26ODfteYmXNno+1jKWd85D5cnJg0PFTVqOAecIPqXBLtXvzGovq5VU67Ip
nYSFyX48EO/GqKfnmOTCCPIXxwhu1nlKkUJ6JSskKBsf628RPcMCv6pHXgY/SOHN
Jrq0W+EclqfQZmJvHQCBfRNyfE5JSHmBcZY8MDvvk9S0Z5nd6d2+b4Wq2CQQcze6
6v77uouugWrcpCLgw1AofDujlAKKvXfsA6IVGJ05BbKGkNN5CmK66HcbS6xSgJHx
cua4iaG45tfgrNRirgStw9UJYxGsl8Jn4Ax7j8uZUborrelR/Clqx2Y2tg4MO3DJ
BCYleHHE4beMCB/kSPXQjDDMibGVRq1ZuQ+/zd6icaUD0cGhQaZ7X5Vjatwbm3+m
LAmLppBafsW5IaiqnPOIZnBFR55gv5H+Ks4J5OzMmmk4mzkt1tshNirTO2WaBcd3
ln5hc7IubryunIW3DwzJ4gcoSLLwgeqvQmCydv79fQx17fhykS1KyFvQI1GEG7cS
DUKwHRC9S8KymryLshiOK0shpb+91nQ28flCBXWrfHSbJBwz+4QvoakRaCAwaoQt
xi+N8CPuVpffU9DCKQmnKzQ7EEc8rcA35OgMFhDcrENK20VoI06xvTLf0ncM8Ynu
Uy6dnOXFEQ+KQiTY1xaaq6TF9g1F+bT9PmjsgLfBnCupOBi0mXSxZA9T3icxcp7a
8HndKwrUUKO2GIa++UWgj5wVKqpxYkEtDQB8XFQNl1XcXd6jLKlT/LBCzgilXRuK
rmdebNQtXIUMPs6QIgZwNHyXPHJglqFa5IsP553L5Kd7jctQj9eqKG+nzGwai5rY
mlmydeBV/z4shKg4OTzJAvwL//jYUktKeUpu1rY2LjHGCuxjTPawTopnnnR9tXNI
oAszVGtjJr5M1VsW0dJHlL0GuHMiqoDDHQrdquA4MvR3M3kEZH7aLTGsmGUylC0Y
NAWn3Zc01ouq7AYz+lAeQLFQ/Oi+piUtXEtsvtYCV17nsW36M3RdnmskqDJhgDYl
TFxEZvhTXdPUzUQZsX3CRdusiLHXqwEh6IuS/toTEcHzvZh1gvbgGI9yD/+OcJPe
f2inoLSsoewhLAaXqMEv/IjF/KqFwWUFUSUl/YqYmA0qj7cZq37Q6DWOzlLy/kLI
Zb2ztJujMHJHZ0AA2jwcPUatGqjlkFexnNd4+BhdXQCabok7LYBqJcDqx5wxalzL
CkDThylnb6UKM6FQabeFjzJJGltLJlW8aPnQhVey7L5cWZk2/d0tbjlBcRC0+W2B
gW44+xbtG+aqjZIU7/wYBpae2wkxI9Dzq6ADd6iHXerKHRM2tV1UayWxZY/XaXvg
b7tmM/n1oW2Z5ikxqW10pGnkYjHSAQwwV2H8BgRYRaRPu41BSNhHugmIFxrzCoTW
h6biU4Q+3R6rjxtvpDW0O6W0nuWrDDLRyiXg38CiZIBB5mnlFZ/TxdnHN06wrjMu
rCGxyNmfEBXPeaBH2HH/necgVh4PIstDAKKFiQP9t06U37F03p3SZycmUlJQsmrt
tmWr0Ls7q8gI8ssHk37N/XqA8DGurPDYEj1Bo2EUzi5tG9jG/oljorWpuiK9ctFC
/pgwYBqN0RHakXLtGRA9AwK+Qat5H0YwVkzNDLx8wPlyn1npKG3PBXaV1VJXWtUd
sxLso16AEgrhJmhEecQ/DZ7Eslkl9BrC399M9Ge0yFZr25GXC3Wn9LupzI5GPswL
DYcc1MmaUrXgi2S6LghOliJHa0jxX0LbZOrgLIpuKF+EdiYCN6QMECmKiC2dJEZF
3Q2Ip6YmsGzs1G42syZBfiQlGTo9oWnjgGmNH/4mOIqKIv4Y/bHx7gbdHsLvXaJV
DmP2gYEKH7PkV1TRXJgXSD90fxFh4wMULEDbY0inr30NV7itfhlaHF/DaWDTkXhs
9YdvTq6SP1M1tRTibgcDbLUATy2Rg0OEc6JW+LjYvr/kFn6qgKpSrEuGym3E5aKy
z6jbMleOvVre+/+Ym0rKq9qjbC2++NOwKu/7E6GWlFdSyWVFx8Bkncn1iSKJ4Z8U
4fGAFekwjxvUiauHCs1VgIE2etVP33Q6opfdyNpX46JiS9JJAXAldvI2vDIzGz/m
OG8HkFvVsPYWlETttDNOgiZ1uFpjNkpoxjU8CfpHRNMXbGDUFppS9MPs2CLPmKX/
soW6uDU1WkFHmH/iWH9CheYO3Evjjv5c1cRc0xvfUqHuc6Qucq/4kRRnVAl5Niyx
XEvKkIFTeek5Xq1PKmCjNKqtK9jbrHedBEkrfBSPA+jj5EI4eXXjHKHDHHWLErOT
VAFzg9+zogl6osclgVgQTe9zwYeLxNH5s9PqigncBUWGwEMCBmh7N9Zoau4Qu5oZ
lTNmsC5qooCn6eGgTfr1+/IpQmNffkjYMnwRNtREHLr0TPVrbrp6/kP+PfT5qh6r
ScmqS/J9lopKobZJGFpIQm0PSm/hpFuCTWRxJH2xxEQz3u9/+F1VwDT5cFXfxlCP
JeENFGjKx6QBsrQebPDnsHhKBBDG86gt34bZG4vIVvuhllgZ6JQIeLkEULCOdN16
er+uNrzkMTRrh+ZJBZPVeRvzl5dRy+90Uleq6zhgjTWXwoGXhBJJ0DrFXTHoZDP6
ltjyDHkFyihB295MRk5K9ver2P9nfEU60Jgw1hJgnzmnImvFjJ+tJ+uCqNdT6xBQ
SEA7Ptxe/l94HVJtxcA2gTvj4O1mI54erdEFUOdntxeOFoyuMNbfNOe3lpFVFj/n
aD1Edo1DBJ0DDdlJUfTHRlxX5uqt4X5gjBdov+Hy0ArhMQNWGlpoGbqRwA/aURlj
7QBT/mBWRv8cIjIMmC98smoZUA+HT/4K9D2ZMI8YpxvTA1skXzSabCFM5yjb7pRK
DmV20mWME5q8PDIqKhFqKtTTycVYFRhR7BF2g/6o+3LhL2+FIBp2EQRENHMtvjy7
JyMuhjAUbqv+J1jc4NXgC2z5du62q9jeFCBMuiuTU5HjLX2BEjN5VKKR0KlMuoy/
C02V5+XlMlYmNVfTflxNrKVYgbcjxpR5XwGlUCjzsYckGs7SYS9+5mTVehG18iu/
Ye98QXrwdxu8BTbGWXZ3WWUYPfQ/Jt5eXRz2m6UQJBCQGqteeYFjK74EGFKUXtdG
CIqApgx38wrRkwd940nh9JyaRmZY4NW+o5wGTtn9Bie4cj6zgTEY7ftmhMTgL3j5
79qj85uZXzF9nS8NXlHE4m2m2cMZ/n3JMAPHxplXYSKmt51w8q7wh5mY96wcbjwX
F/DUm4gLMYRo8ywULXbapGSHLS5j6RTzG8IpKbyP1bC2rvRpAvESM1xE42qz8qyB
ZnkcTf7aU5A3vKDk59N7BK1XRwB8rustkfeqs1lMVd2PGErLLI2LmbmmuCqOjeaw
3jxRWOYDOLuURedVmTZTyIS7n5M78JQbECwJoR+DlKGPOB9fBQfJ9gv4jE2NFGTs
P1rT9JK/k+BrpwUVBu7F9m2tiuU1kFKBwAxM0HuVenJ/vo8gOjghr6E/epKkHblL
u4aqyXYYisG2JzmMeCju0UC2VJDCM2lDwIfqL6L0hP0guuuJppJpyX2yDsI5IAfo
bRG7GNnYBUUNdLoMOxtdg4t0TgbGIU2XzoE3IahAn8SW8JYH3f5jcTwAxFtWsDY5
x2Kq5s9luIva6yRz86f1VV5efbibuz/31SGslwWNUdqlj2+BzuvKsqc93WMKtq9D
TZBXmQV99W/opzcbGQxQFTJrLaa1eIAacVvmNneOTZbZ8RhN56GRz8Ze/QbfLzaB
W+fWCCP76uMrKkSRWb+HUa5MJbKJDfnTXu0WICSKpkae6HUoC451JJFQXo169RBa
Ol6ovKGJHIjJJqRTZBVwWbrO+hw0bais6CLU9fbDFRv8DWWLu/7eCK1ffJLt189V
8+sXMI7Uwgom4A1/HgGKHGS0jkT0xfzMJ/9IquNadefbcnrZig+ogWQ0PSbf+FD/
cvQ+BuU7sGRWGk6N1asIdmOJOXInoySDPLDBwp3MsDXlB/RMsLpoVlRCmYtBwFox
eroesI2ulIvYTlpvuZrlcxwA3LkBAxdjCAQXZhWF+sar9Q6wyvhfeArWW5w9Sjz8
1lI8fe44b8FqQHS5KgMY1SRACclvqyyJiPbwoJj/WxKIqtC5RdT38LsQUEkdMtxX
MiiyasMVfyX/mpNmyUA46XyUUKCzD9HPCLqG5bkvFdkXS2cSlBk4YwjDzdPJGBAY
7lRrHTtXh9kFP6UpeXJ75VNCPKnD6lA1my1E1wAAf9+E5qo88VXZfCRmMmlHuLqC
rCUK3e3iUt2fleXKVci1IJbjHZ3UH0jGJmZipxX35yEIImhaw0StMc5tT4PvR+vC
ND2RurGi6+DvKSYIhB/FESZZf36D3g/FjMnV4LZ0yiCY/YWKw9clXCtfQpyWyevr
plwHte8CgXqiQmdHyhcLVgGkOstBPUbHZJD4hgbqFiFSIBSj/dw88p1cviL3Zr1A
7vLaj5AtOdYQbjTXPlWCzmMtnIpw1ZNtAC9TqyGXIMO1gGh/nQpgI1tcIis9uK6C
NTbCBQPGX0YIBSyWC/TvL+9cQvBK3gYfLaE/1CubCdtWWVl2UHC2G48/CtYkn1YY
kXHw9yCvZ8gZcn0GRBYXnHGftBWwWExA6VJB4o/wzJ0FMu0Slw4aJ4nHmKR2cjyJ
AgK8b1CfUUTuwrVYT4e5mbisbhmmKjpKcEAemoYBXsOqF5CImHQINcwEbg/0vbDF
tJ1C3spGgxlOxbTXulFy2H8npbTYuU7q/0MtWDfK3o/77JD6YqTMhlmM4aVJAwX1
p1l1a3SnxsXqunQrcR0440d/GEYgcxwIvrtzCzmbIv4Kn9ZTT/C0x/0uMWpWtHX1
9PmvG/hqwixUqKr3r2Vw/l0KfDQok74bwhgmj5R7qK9/+TmwSkJhhhPHqipY81Th
GKMEH0l7NeQRqci30mqQhsQLT8DF45JHtY73TCxnOFFytA2iQq0MzgFa8m15pQcO
x2IlZS5GaW1AohN3fuaSen/p7mCSjOM1loJfpAcVoN8umyd9Ng++PJtoOpnrWYJt
93/l0X6nydycbOMimmBh8uLT2GujQkHaEK1WPLgxgtCoaaGTAeR3f3zU4tx+K7Xi
gTDVhuJFxl/9zJNjhTIwVHNcd4kqMFLp7KC8L1sYC9x/qqTf3FN1oz1his+oFmK2
pO++rYIYBr+6zU5LdAoacokA8tYMdfGG+DmP/3qt8LaDlRHWzSv35ZeEgPRI9n2+
KJhSVoYxICqAYiUl2IQ/LxkJ+zyhElmaRFctVGC7qMmC0PPn0DXpw6Q6vqHGj3cW
zUHppk7EMEzyw9nJJr/7crCE6S2TZeQGbujywYf4EP3giKO1eKhY0acgvS67SlVL
InP8VUfNWqYxZtUpySEQn1mbmzU6enCcYqT9mK6VdnPSJX/cn0XM8oOPpa9lrlaU
+0U7x78ud3wYR9kWVhK8f+C8PqY4e6sAIrDwbPrp5zOBjS+5+IYu05B2EpPi57c+
0wtea9rgBRy445avz4O2M7OMPkh+8slocOIpOclgFYYSYLtiJGWe+IATzrfl4V3e
JPJxzVqY2MkIZff3D4Uww5jS6/XdovKJfx0EPJc4H3nbvDC7BX6bbBoSA2vd7Uhy
/mbRgIxySJeTw+sV1V7GCOzDh0PgmuV3NJtbEe6jKBP1ZqUccaAm9N7I5ODfDTb2
4uu9eLvJ7p2QhbAoLXM9N0SFwrnNjGha6AEH0mwXg+zIuDY4A+FSQ/JI+iEF0tU4
WtarCiyLu4IG+zk9pWfJ/ZBXvDNReMcXnrq9mfGNwXx1F1SoSOYz87oBL7QOYZBY
77d56KVpve6Dp2xeEYYDnELI8riZ3IG/J6ogmZVTv6M0Pnq+z8LIbQG2CPernHEz
xvNs3Qx+jpyyVh4npMqWB8o1EUK9E2R7mSCqJJfqjgQKtq/7tYfO2pPqfaQGmc64
0ZbULKbDpTJCb70wE5EDDAQmUe0KMe2uwxG4VUAjRqRF3b+/EEbqzw2TMgY+hfN6
i52seZIlw+HnFEMfj47C4ZFq+rFr5KchQNa8y/t7Pbu/2/ItA43CziMPDhjL+aWA
O/wVDzOM9rDoC6YRfqSnD512NixtgvC+Qbw95Kg+mQyQ5j7ZAaw0+KpgJpredbpl
dpuSnO0HxD6bJiL5LsIS7poU158xw4jTfARnIIrdz5J59ca9yQaYUk7ivsUzRP0B
BBm5721wxg2EkuAZpkgvgOH2lOV++X6gwRNxgWCwhzIwuD2DT9usTNwRM8aWI7CN
JdEckK7URYZxgLa/gEjtqNyWrSjpXcLovnr0fAMbBVPOzEt/0jWsWgMV3hKC7osi
Cj18cpGHUpXaKRMaKFbwgTg5iNbs51VOXxf1cosuJh3J/YO+z/OSyuFR+OpJ57sA
gxOu/Y7/OKZPIM7tK6UzNoPGQsjrbe17aw07UNp93GfRIIb0gHwAe4QJEWx9AEv8
qecNyYXiKk3qMvnzbEr9yBlsy5drqkXYLcQtsnK9x3IWawhAATszGs59N8arwnkR
En2siYhE6lv9O7Lib8gX/wmQfRhVBjjwHHC4Lybn7ZBfZxW+dZOCQ6ajJAyqCJCv
J6r6UHWtPpv09h+GYP+5RMaYsJW9adWzdX1MazBtEC3YLDI2eoC5QX7SwJUoLUiU
db04BAPpuTtecjIuPKoL3YfG8DxHrdS0canj+n4PophSxGRIlU6EkTlP4z08rdsC
HPvlAqMWs/fprGQ4Svkstw6Y+UNSBjbZm3b03qXkgMSYRZx/neL0HUR28qKB1Aen
gpbr1rAR2s1MVtWwJm92KXQOoR4p6AnbLpS3ZKp7Ya2PK0JHdfwC+PVJ7x4nblE8
rCLigJJU1CHCSKDTvZlkX3XJm3eHtuLqt1D84whhMEbMU1x90jGC7ic0wWRiFVjC
Qb47NXuVsP4o0sbxaqyWyikmoPBIu5JZs0oNZXkMzwSCBkLiRzNbTtDgwIknV2E9
MRY5iyqNd9nMA3UxyZyapGlAQS8gYVvx6NPesT/Ysxjx8tFKCQptZQimTP3rv3hp
w5+d2Wm70DOht2mBV1GvysKlzaKEjlbcw833nZVNSWZCuBWs1aqYEQp2PxqH9Ozw
`pragma protect end_protected
