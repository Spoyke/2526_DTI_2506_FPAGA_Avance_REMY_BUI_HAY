`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XBOjRkQtDa2me4R44X7edYTe9nZucChvvtip2MNk8MJPIwtWrRf3g7kE0qoKPzIz
aKMaPSKoA68Sj6Tq4DM2tArHCMub7BzZC1bGxM3K1KCZFgb/H/KlEYRj2ka6oPQW
BA9phjhR46yfSPWnDsSL+ThrDopID+6TppeIaQzjrQM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37920)
imSOa3zEMD8IonBhrZQVTwoVcEq+dUNNARdvLVDtsYqTPJ5tBKfPQkiJ6HsjI7yq
2yQi8gNddzameNmvoIeY2n9dFD3Cw+DLWR3t589gQL9Qa9f97BDR6mTSVlfkO9so
KhvaYa5dRgTPxvWwc8t0kKzFmN6lZSsT7tZD0vrJoBlftuw17UNQDRuL21VwQAH/
2/Ykm49v+6O4JCDJHr6eXsBchjxI2V29Slhw+VOY2sbQft1hWxFQtlaT8+TwcQKg
IoK5qwFaDjJiRGeNIuE4zagBFyRhB13mKGPap5QwUmxQahwmynfp81UWWUC6CaDN
t0sGatNnj3TOjB+997h2O4epxffNrsdW5GV+9nIw5FovOjfzOI4D29nGkgAcTheX
Pt1w75vNK4Lpdx5G0S7YruOgD6CxACUL2AFvERo147P2j//he2RBe3gX7jtVLGgu
epyEGahClHRe4lDKnrNbSqqYqDByiBM0fWyv24jxQZy9qXNZs0rJK26IoWRoBFEw
36oa3kw4fox/6KpRXZos4EW3TOEA7xlM6fxgRLGpQiLF3KIzFDXCRi1GhcQEyQ5T
q4P50MtYAsYTGORWRDeyBk382K+y/MqEWjMF4IG13zgnr7ccnp0VVhRFCFmvRMvm
c8Ls0FhsFeOjOcVaJsg0zcK6UgHeu6pTSNABFRdrbipGTFvfQdWhIdgiNjbcLqPl
UWW+lOa8lPlxBOWfl3dr5xm/h9r4LQ/MidZX8AzDWf78JXu4xpcBz+GbWFAEkoV9
GfwN3KmPqnfoND94SfElmrbDM7Mn5U9IZa5h834FqkwqZrqUrEFfyVf56B4DyXv4
nbg2QDXhsFx1tW7da1+K7ohixwyd6GFXpKc8qagdsovqbPwzkNiWzE9hYllBqI5I
KnAZvTjj5sbtOZQyRj+dRhZ+zPTwjdVU1jB8ueN712eDW/23hdXCezhSwBXZbjEf
oDfp17rbewroz2M1Lb57+YFmJrzVhAdpAI0YxqrPVUakdij7F1JneFYkhu2EOEzP
M9DMlZTx421CSsBd5BUZIeTKsRCoOoL+IdtFm2UHSEOC3CI2lMj24locdPm86SW0
6M2CiK51jy5tEXGFS1IRP7YOAqq1//6WyfMohAhl2a32/6byCjTA0cDmfqMSXuT0
xyxdUEuD7pKCbLIwnX435ypk/V5/UEaY6ZEqs23jXqV0KVpgnB7/uIYxUGbEbuQI
wdWMr1OJIYg2qwnR0xGjI1n3384w2pY9Ac4w+Vb8XhDBLrfj9yw0u6yKm/ev8FBa
InZdj40PFMJU+poDWtXawhiYeRqpAbI5ZUA8ExcwjkUbRcZF+sGemnnHYy44Pgz9
QQO4s/0dPFn5uU4o0ifvBoo9a4AIIK/Uf9J+RLYYhczwDt1vrSLOcyfwvHpypw2P
kEenY81+ZGyQ5NsynuK6thG6ODYR7l/J1I6cYYiQdDCtwLOEyhO2ltOLTKTMl2I9
aRgwJITQ7A6mLSIkYE4TWeCnChwGW3vi/BvhIOnH7NkqNhv5y1cdiZGHvmT1gZEU
qI18jRHFyqwT7G6Dkz2L8K9T78rj1EsXMrknbWtiWjKXVamBN452ulBeGWjkWBdQ
GWTQKJF9HilHRQlMeVpIaBSKrwy9M4W2Qe5IUUVXy5/UliVuAAawh54Kszho+zGn
FoAWgphkDfXegFU5gz4CTRMoOnkQ0Jk3qKvzAJdHeK102Yr4Z7vseAiHH8FnMvsD
tB2szjZGBPPQs+MR0CP0q+n2Zu0PWbXnfkmN3n8YeNP+XsGio3jqcqe0ZwTkUGi4
lmu4dg1/oRBMhjelKXWIx8cfB4xU7cFeYIbAMY0yYVkBqgGd+9uwlhN263xICiW4
Llh4WXRRyZgy4Jcippj0pv/x3z5TxQ0ttT5X7iLuaGLvxPEnU7M+6NK1gPratdYW
T8wusjot8f+ezKwFUHTl/mfrHbg3B9aq5frzId9Er7P06+gT6ounCkcXb6G1N5lY
bATU6Vt0yJFY3O2ukW7Zza4TVIfgCKbEVezY2DSGcJpTBkDeXCbfG4vnUYcGuI/c
p0YO6QWBq+Aeiq3ZxVrIvgQWh9PbW1GqKA+DSIEYfiDOEWOgMEI/8AvljWmbTVe1
p3ZlWaExl5Mm/ogNaD6HqgC3BA+TtPLsTCK4bpSdB2MO3fqDCCysMpCnBWfMW4bW
x1Tzs11rR0hdp+mB0ZfGazFQLII5rbyjo1VgvdTrLY11Bov3M/lDJ58ywMIYog4b
gz1OlKwqrT+5jGc29VMz6a7IBO8gG5z6++DPOwMdyuiKrAEAMNcvR8JtX+kbi0bG
etPFyYURStBmI8plR3++EHqqttauhp1gwVa9UgcJuuQJ4Zyl/jz8/vVSvYTfMxJ9
wsy+kVd4+CDsyKq517h2k4TUHEYHxRGSnZphwg3Bpg+Ped64tmaynEj0L8FuDe0H
kJhqucMYes77itUyysvtpi/PhtCvB7+5PBt+8x7E2jsIRYMp3u/MbCs/dhpUaBm7
DeME8n9U5+axBMGTSm1pREGpBBD0NkEkBkXNPI+u6hrp8baDJ4qX0/aBw4Y/5qh8
ylgCI3DGxNyFqWIzCp5byHCjlX0jMmewsr77x/1VnBhoCj1+OvjWD5xv5XqkeZ8E
ieTFwWAV0L/2HNsbhJdgwCEsq8gqiV5izOnFolANkZt/vHz2VTgjuwmcnHMZV+6R
pDSn3doUTfJf0BhLE2VPgbe7XdW+sKzPWIubGozDm3B65qsYHTafizpKvMEgNBeu
s1Ujs6L2JXqu8gKKuRyvQL4fGxzUSs/ZDpdrA0cxZekeIEkf/hTnAMa/fKQkpHUV
QbVwURataOUKayPjpx3Yokc6bMMV1vQ26daPDQy8WsBKwyyjZxn2j9MEGyQYJY3F
ZtGPvpuonulkkRXq1v7Fc7YkTw3gLq/wkf95OfE2kPMrF1wSrXDH9CvHK57JK+OX
2e+GkNxjyNqIuLNvuAw4P3xKGZRi/Jggm8pl1k9qOTRQnKVKTSTwthRs2dErWG0u
EqAAuLAbdFLaH4HLoMFKSNi9TXl8TiKKes/Swj8AshecjmjjaSOkmQeHe1mkRKE5
Q46H/aEjAZAF3BaMb0M3J+n89jKtMZ7UfMxCyPTGmFHIm/arPuxT+G44ir2StHV3
vEKsIwDQbcClCv9ehp1r2e2gxnj0dalkCpbOzetUNNAhNEcW+ZUCpzYnDGuljtXU
x8zf4rHrQ4KS+aamYyq7RQvTf5qcI5PnyElbzhidnqHE2nwsVzyLteslS5S6C+2k
NLzkvXnmTb/2YEOm5zyfzMW/87Rhg1oFmPnexGsyEPLjopoMc9a7tIG6EiTwSoa4
2iUt90oPcB/uZqmFCojAG01G9g3LrkqkyCCvQtllNvK0yAU8EVJSYt0lUOxqDwxY
1XpvQkCe41G8TaWxMbXpSxD5wVY2R6UaXXBe0RT0UrAfQ4rc3MTp54WIJJECJSxA
/mKQ0dCvus7O1B1U4nUgIXl+yNqCCEqEZQI6pZzQPCGpnZEZIFJIVI+kf9u7BUwu
YFQvr1utKKU4C8gaX2jXGWvX3bjKmMaek0m+IcgoeB01lCA+pCfxAbC9bM9O0i14
HqReGLk7+kx91aqWYHt425WB9kdbwOy6pnE1QiyGqjt69wHO0EGQKP4fK1AFYneR
GmDQwueXHww9ZRBEeJHyAUIyzk2sYPQ1zV5b2gM7gBnna6MNtRsMd8eLQbWhxk3S
iXy2G9PnQD3N9xGbTsqMYOrsnOFEZe0dkKLtdtiMAMEYz80gZuK3R582GoiWMJUp
gfvW5xW82eZwpp8LcOF8RH5+MB3pA00jL73E+ufmKoLhqYhfJ/R4GL60iRDqSpwY
pVFZbgQD17sdtYYhAtvVEh3ql7q0+/e0TEnkc41LDfQvJMAkCeBJ6oCx3TUI0hFs
L7km95w+rH5oUKvQZkxMu4zrSmwz9p86dgGgOcsKga1oXRBkmU2mxF0HFqtqen11
EjR/7BITR+JBDRK6wTP+2UYvk4lkvixcWAVk4+sO7mZ6+wgMsQh5iEosujKRSrta
At7qcbo78iBIATL6i6jdkpGu1eVGPExK4VjHByANqbwFbRdRztu/y7MwIFWsB7XA
+dzp4aFX+LseLjh0O/PJFT7eVeQd7hTB4vj7+YwqTnPJauMQWoJeNDK6CV7chjEH
ehvDn6nkPNwFFfr2T27g4yB79SiBdasTr+S4BQLCD02jqEE3f6d9HrurEzpX3DQQ
LUwn9ZWmlwFSqIpJNCnFVKsFc3xMmwX9EpW4w6IG7pyoAI1UlTvSEk18Had620Lw
UfmnKEQEYKJ8navnbxXXopIcUlq/yISQuD8VmZp84zuiKYqSubXDMV2cjdbm+Lal
O7IQhJ/eXXMOOGfCQIV572R4uerkXTIZ8Z6k4qX8hp8zdKV29zbHQ5h1Wmoj9TYA
G0HsxVkASNFxebTVcUKwHlu5uBFgghJKytgYFrtD0lydbVF8jQg+Q+ACcxDls3E3
Gkvjdh+Cyw5kRL2a1zLntlG7AHUbWcyMoNWHk0I4Ayoi4FFi9154Wp9KEzCZHeI3
OVoddAjRtj8Fj7BGZFlSv6NZ8bKo+/TW5aCg6hS8skt+jxK+NYqUI0sNaVAfhPyJ
/gz/dN40uMC9j8gjPWeHc9wx/NkOAR1QzDjwHjEIBt/FwhE2m+50tzDxqi6mI4Z4
E5hjlM1KlteI355k61NLx/E8UTxgjQnY6i5EoMfXjzWizrhXckD0iTIaX4pzgZdD
LrTqaqW5DviKjCJsZX5Knh2+SU159jwx46l1+qvKxqSmHist9uOVbzZf5c30iIPI
6LxIBlnFx9qkNWDlVW56jlAa3KmYhOTUc9XrvPKhRlXClrYlyNp2y8mC0BheUJme
FIdUyB5MTplS5wFpFmHsBLY+Zq+0FFNmuLiBfjDKX6eKbkj0bI6ig1p3YgrDhfkQ
tAX0UPY2+XnGZJ5Q0TVXB+93lGmKzjn2iIup3lVrvU72XG5LdCCoHJMjt7fOR59a
yK8IcoMEzdTXGo/YW/NpvpJlDqEcQUFW/uHbQVZ1ORwOIhRNL8UqEHRrZjnU//Xh
abWpDZ+40JxCSztGq40u1d8uhxNTVIy3mH98OvxWuKT7Lz3LxiugdXbL6+GFrubY
D+FkT6mrAXRIENwlCwU++KNkPk5YrSiOMny+Bxgxnx49tj1ng5DuUs+uSSzOYPFy
YwRvuNuCE2FNyPpKNUwJXSYZb93Q2EAGTJWaHSmuNHqwbs2L8QvNCEX8sbjRgIfe
GSy1jaeA6F4Uh0oYZ2EsGAqgThTIsSETINXtlGuCdRw8q0X8LR/HgI8hLfVmOsec
CTTH0n/vYkM7/M0TodDCG+QnyqeubPzQMn9FhNKrWReZYVzRi2774w/Fm6iuzUm9
KkvdK7rMxpRDgQBsNU14DBVSfJzbgD1z2SOKobgd1ZIYfLeQadsf8nMIVPNbIzdd
uVV31052APeoxsvyQ6EP4QRMlhAT3DyJt0t4W6Ju1o2FvCHCj4uPivEK3QiiYHw9
TtRhlrphRtH2dygwH/bPKEpS51iI4fx8SJHCyIR7nOeplncpPrQXCaUKm7rRnoT1
Lb3lnSHWnYE+1Fu1X3bH545h9ILGXbVfoQ6rkaJUh1CIEm0oGDm2p4B+R0OMYmmF
VSY2FbQUA67r6SQCZhU19I4WX7a4qsuU2AD/D/zO4PX9q7v13FsMAGyBw1rJxybd
A5CcEPCiYk20VzyavNGngCrBbH7fSGlO1y1hy/6ACUjPLKx41DF336ACve8d/ii/
QaxsVPJA3FyZuxzQOOcYbI46n+/hKNXZlxKrtbi93Tz6XhL0K/wV5Z2i63FtK4kM
7S8Z1ejEEadXOKC1Em/qP2BOgkVjN/V/LuQAuYoDoGpAtqb9ShGiqkeGSry+Tgns
TDlmK5HGETzCa8wV7YDxq/Pg57cz5Q6WI6iZ6+bMKBSi7+sWOC8weUC1/3bvS1Ir
kziHV59DPMlyv+J3gibEWp04InvYUO+2h3VFFROdnzo2DkVzUkwZ0/OjZ0Kg60QN
NHsXMD6kle0eFsXF/jyGp18IEAwQZAxcJynA91loURCCXtdELsexJ0r7s37wn09Q
nxoOwsX9/fEt4swNp2Ns8WMCpQmSurPFHNs0Shi6y7cnMsYG1ByztEAoywMJWe2e
6GN9nSAhgyaEF++/SgMo5tNsY6XwFL+TzPcDzLsPlNSRQssaQMfWkYk+SYVHyyxd
DmYh1/NpoTHV4DHnf5132v3ISKuVclCTgVCX2gsDoiJZ88sufp0UvvmW9xTPxcgF
vz6HaPCRqmHhXm4bUY00KRgHer9qa4ntZ46ZZ3MNiZt64rLOypxzdK0yEY4aJJg7
pEFpuvgwYu0R7QSNRa68N9+9+auEoch7JcWL1TKczEPYhNnd+2y92aL55ML/gpmE
Z6HgAplHaXPf3//2J7EV+APf7BatF86lCR7CMok4IN6FSjaS21hGUx/ZYkA/JEjl
Q3CoqJkbCetV14whFu6KNVPcyG6K3cWuvWNL7aPyJHStCH1NYHuFI4LA8oPCXzFu
IfWPdzOsQD+PQ7on2/bDmyGwjpx970LqBs4hzm/YEDCWH1/Ti/2PgHADHRG/ytJu
75IRXsT4yvFEUuyDGnNZHeOIonTa8YdJKUjp3nUvcgjKdoJS6neve/a0x2kk8D/0
p2jWkNrH5zr6c78gKrS/8sTWumy8LtaHXTqOB8SoqHrMlvTWdVFhTzJcf2RxxJte
dPXayW07hIiQ96dO55Tdf2EKCXpBfbplALRtPbJRcKTPzq1NWdO2Z7S6IRBYV7W3
HldM4X+pYTtp21SSIkBLh7uldgecbrB4+w0mPvNhy3T3gzH4e73wLBp2U92nP+as
t6pi/JVWYCOF7kIK4hhYBJ4Gn9XH3JZxVCl1d0NHXrYX8vyx8USvfidSA5t+FNNk
aUt5Y632BbLosYRmlVMlW1izVnffFj3Injbr3lrxAy21NvKHqaov1xnVJ6ExvfhN
wXMOZLypcmFO7XaPc/YDIodCoqb0IykVwr1NifY0ltSXUHmxYXb4Q9jr5z2pXssm
POb5Ry0PyDlDGmfgzjymVpo0nUlRFJLTiz+Q8qZZYN4HR/YMkA3hEITYACykTowW
m3Yb2iIwbmiO5znmUC3wnmBtzG5s0fxLIWvXBt8apmZuGgDpW/MzhueMyw+eO4JG
BC9Qfvd151IS1WpmFW6OP5jEBg3BGCiL78AN/abhbE39wHcrZFtovpfB179L1qKV
F9IzBhQxFKxGWPxFSiGcXV0bPkS9R1dWHgl5cFH8ezI2yZIm3HcoebPRYxu5jopK
iljkiY98SF1kzMW0IqzFgmqPWgdKkfs3Od5ZiWcxSkCmihCqSj8Howhom2iGjB/d
plTLIp23HVvUZr4VWJCCDpcHGUhye1j/gZmEObQSnm5lVSZc6NcOx9vv/gTW7wVh
7gmklv6kPDziLcDPan2qqyoGUetQell6N0A84xSQyNDBIWzGO4pd5QhLyUuSzK23
JXCIad/KVmHC2mnVQzJja6Q6plWsJsT3lrX9Zzt4dUmDFEBFik+326Hvd8P7Am+/
nJM2miIbOelFNHXEaHvocBWRC2Pa6j0d7GLLuia2bIDGI3B+9MfQuwb/d2Fi2wun
z3/9ZdSJS6FmQU2WzGfjh/WAGkM9R0BSnqwnXu5+oxM3R8RgKa5+tc8AEc2MHomu
ujecVMbn1Zxk26XYTiTiN3NXbxQasbre/kaW9n8hmWqKfbAaISdEzdNAxcPbRvR6
KnoMoHwBgyDzIE3R6iFWufqp+F3VbqedMiSNOFhZkIft39O4rsSVCnTTZK6oMFgS
LNrJ7uRumLkx835KYEmPc5CUCyLv2Y0tDueFUM9d3FYK6BECHNbf7GQdv/f8a8sn
LBKSslpY+a5UPR5QeG3kP5w8LkLpPYzOmf/pOAVxTdZ6u+3yTm6kSFgC7ytueT6K
ClI15l9/mW5d3x1v1aTqcrnSrw6FNwPzZnfJ2jMQ1Gzqn4+pEI8k46Mi3N6lYtdC
MUeDqPUui14KSku4wVRfM2AiyZQpY9Bk8piqRVjbaImehJWK2MHS1EE41u+djy/Y
r2gAjj/kr2x8yrXiQ2PkFzR5iWLEpbdEltvT3joSb51lIu1VdbzSxv64xY/R4/G2
AxttOcoAg5m4jxBlwkQZVkhwHjSnZOP6+Fs0us3iEWhM1Gvy3ciOlXQofUWnEtJN
pVogHRA3OOguSTmhaoPuwE01GER1r+Js80rhN+zRPt/Zmfd6jaAKvwSAcx/gx8I2
YVsJ3sNyjcTQiZ9/l3RssPi5qX6vEWYuxgR/TwuPfTQ4koL3Za3hPWkkScFWQtwN
qFYa4CTR2hkBiXw99OsRewPIQMYAodzeCjzKBsQlMNSyjAAn4qX+9orL1qV8XUIk
y0cmG5XuNBJ7AkLREQ/qdlybZafLB7sBgFP324pBINEdnyh77VSFRj3vIqJxojM1
nPzftfrvuZAP48N+7hRe9LN21Y5guxegeHPdiphHWBLPJ4hncwyK+nK3bjU2IA9v
xwbxm4US94WCRTwNB4h57ar4+biKvuln/7NsxBINxsS1LeVMekKSOZkwOZUlHmkg
TF4KIZGDcFXzO+mMmVass3XSzU5TW60Q3LqH5Sws6fxC+kjucXhXlKvCY+NBTI9i
PTt3vyTp+Domq9kKBUhktYpy/Er4UEWnYdOJbIH4UFO27QuPc7BJD7FvuRwR34ZN
oM0kF5bfwtUE4akXhUs/GR1qZ0rN/ha4TRtZ9HnU0NI9enWNknqGGHWZogfnRTot
HuimMucMbZR8HJZ6s8LDuG0dJvTA3GR2vr7Bk2WAR4e6CGe0iwIAZIWVA4WhdFmR
tjU+gRVHZ0qkcFPkP1OpplecKWMnecRkYyMOfsLpGEcd1U/r5tWd+vLvqqhsjCpW
faKMe8GrJyNP6+O2B0FZzEyI9ZolQiPf1JTljmESi00PPJe4+dYSpbJxjQrtwQhj
NhcSIlnLo8hsjuxbJ09rvqTMmnp6Ttg5ETkLKy4M2zGPf5io0dD/smhC5fy/JVSV
le/QHhWn2o2BIs0f+RK0EMMac3bseFrdrFLnBlIfcOwBWkM09CGrwFHAZNq33Ouw
+GPe9ESM97H6xfRhbECykijm8oyNVmqYmFMLbEbAHt+/R2Y65mEzPQQGn6HSnMyk
bp76PKNN30sN22vAzcIF+HB6+s25n2ThXVbFFArqevbTcNlNQlyMc6QMhZYEX99X
NEuCSi4jkie0a7oYo1a4jbFU3VbCs4UQIpbeiaGmY/oJJBBRA1IpobmGwyoSQndT
EMANzGFiy/EAHLgOZMJYk3Yba28mHGpUPdjeMT8acC3eqs53ASRASUJBzg+IRYwU
880AIe7DmzGO2J3t1JpZvckU6wGUawvf2tDdxhaRSugGg/r+XtrWEeScstvzVkMr
KjI75cJ86Prcl8MQNr1F+L9ty70CtQ7k0ieWkFPEObvswUmDyqqjT/QJMWISHGqN
tb2wpWOFAMkakYU1aysWeMQLhgrXzdhhsK8blfSGFijTxTWMlYhT2mgMkfI+UlAg
AreSgn+M7wmQt97dprpKV5dP9rkJCSOGk6dzHemAzM9CGi5jqQcYqbrACmso2FVX
mw4ryLTo3yFB8p1Pa3sm1j69mo4aqaTB8alY4cawZ7midJPC0kNc0knUwDgyYjMG
vTf1ngVEWFAtRFCivCL+xDlIhzl7c4FyAKkeo6YSHRLBzDRmoZcfElOEZkpcJwuP
FIccDspab9Vq31/ga3eIwyAMV25S0C28+O/t94HNY4xAk6GzCSW3Q1h0ef0vdj1s
uQ6k1o52vySShhJaJm2pqaRl1LusljuEchSBd2VWeRj3aVLmsTojvw1nTT2Mz7ee
b2hbqwuWJWD7WNyhLaG6Hz3SDxt8YHKhMmaDA32/ErFKhxXTx+nMDkNJ7xaskRq0
vLv2XY209UN3kE//oKydSzna/FRz7Bv0bhSuGlyNmEuQPqCm946JB1SdIyVLycCG
X1U08E3Q6G7ld9OM4/QQo2LL0ahh6tzZNJQ+NP5Wsbj4bwy6XxCdqnb/tJV2Lk3j
7PjPM1r9XHG+1zqZBZS/Nx5PSvQfi3Y3hblLHLWdXomjUNN1aehMiAote+PYpPJp
kDlWlAOk2ezl34D1covmwF69z6af35iUn9Q8YBG5TLZwHVuL1Hzn6ADDSqmyTu0H
FDFd0jTMT2MYJTSy5VSsI6hrTw8gHeMtTdAvucahqmIh97p4tYhe0Go2GoYRv9oS
sjvzsOcOBsjpVF/vYAE7eUk+JLSUp89L7MBdiN3ntmoB0hm6mfhNyP3QVhaXXw54
BHMsG+EG3TqKTxDqNdI+zHdxifDNoLTxQKfnLYWS9rrgbb1MSdO8sGa7edKl5Ecu
l/x+bzGjgXUUzimhVy3sBVPhFOIByifsgEhbc9wrJIv2BuHtDDA8fiZmmu7VD8Xf
SImGyZ2/tw+cycixJOkaQbiUNuvlhq+l76hsmdTZZ0vD6DL8MXOFretyWNQCOJ2P
b+wAkU6TKEgrXsZDtjKs75X3CcdpQEQblwrF0iwRYp6fNN7m7RmbkvTx1BzWWyQh
TC4fliv6Zqa98yNGIipKUv+fpVeSGR2Zqyu0f9MVMHIgNddVuwkCdtWeUBkWOVSc
Q50NbPFMqnMxQTS8VRkJ0l37HJcI5LdNzD0LZZ+dv7BlTe3XyfCom8KSNZz7jvEp
badBrh6hYWu2KgW1LhjCEXdJNaDajSp2tpU+0WVbI9OSs2WZTujzLkNHA1HDY1Sm
RvqZM4bwRqR8LVpvywyA40u1BtpzGkqOApZcT30nF/7qH5kCi1vqX2kTee8icbyZ
pQPU3nBnMuJcvxPPEcDibSZZsR/p8ek6Ya+fAyRwTEloAHphJjO2iOAy0ae0veLV
vEB7GUAS+ZKcOdHn1OUVA6hs6ig2aSGbEl2sewgf0A6F2OuSeosKqMuKguhci8G7
fMSO9zyMunoSk/Zlk/VerGUciSzERTAaHCBJEWEYj4/oqoIewNLdVGcmnkHV5fR1
5AzL1O4ZQErhacgewk5ZXPiQQPL+1vvdUQChh1D3wLSiO6W6l4COxhXOonODCohl
kdU2KmJp1TiTe8wajYgEtUJA57bSE7Nbj4E2YSmAsTusEx5NuxUikw4HWlZrNelR
q4U4Fr6QimihZDkVrrBTiDBLMoxW584b5rlHk8E+VbYZNn/rcafQnWWDtsTaxdYo
xJnnCdrcfDEgV9Vq5Mf8HzgNxTjLJ/22RoZLKwdvVXU4PPJNtoj/cx3WjnPjsnGN
NwWab/PK5xRZ/+ZwHAISXspVRO5AE55r0clL1Lh2xefs76Rpkn1zMM9qGxSuwgEA
CsFQEh7hM6oGFXV8htUxhKtT1qOv0BzbBGUosVp+Wv+7xOGmLWc8Jh56IYwTEVE1
DW9rR7mIvVTMf2hTW59Jbjlx+FAEC+C7XhOezl5biHtxl/BCVEKCch3fk99JHSPq
EKJ4elWVGPihIQ2QmHuzM4ZJqYVS1Qt0d7jUnU2XHujN2duz9eeogVbD2+N77/lr
hBLWD9HNE3R2NIFH3uhBGFeYkCJAYM6lUICBEfaXd0QunBNrk/bAH/CfDT4usT40
FVPBIjnJobxJrAJ+gBY2zXgdTALiYRUJOLmPWur3tRa/YUxaWmLTNotX3xJQuZWD
LmdpYyahN9a+nN9J1ydzpsdtnUTfcs9kbFr+RRTKFkMFkMH2zztPNOPVQBoyZG0m
KKvVKp/+fonxaQ7nKD8A0XzDiLrXKwlmNEjjk0ZlegIXhyjJPpl+Z73qZh/YQD+z
wLf0ncSeYlqTifFZ574c1Zkwm3uqiIjZdPCan75DLYQ7YVMGwjUDfGHFSSJLZddB
/zUGWthcJ+4NKsr3gRZOeCJPwcpdkNdaJxio4dg3DitBDgfyriv90Hi6JvhsLPKk
HfnbjkQ8czSgGh0NKo28THPPsWGXSMkPPsGbA3dtzKqH/iPm8/qp7Dc7LVgVCi5K
8l2HDb6H++eIx/tjV63dm6qt28czuPnmlMFacEsBpv7XI5FuU/JXSZldEaIAi/O+
OAvpZ7l5Mp7XqnNB/xl5KIfbKT44Ms9ncMv81q8NbINtotQCprzPE12yjDfuDoFq
ZOVD4jKcX4ciz/yXxM45Fbwr/EWtD9Kw9/QO6grC3AUWOInuP/345gC12Gao4zCF
evhvM0oF0wx4/QbOgeOno77+7mGuz27nx5R78QoXb/T2Bmo4/kpzBtxc7ZkTgP3Q
ms8mDNf7CNteKwFxR3X/Yrtx9G+bDz0FwryHOTEhtZk6mdMfMJTvPogU4dlUcNXq
VPd9/Dy0BnWM9B5wgwnhPYAeA+JFMEhz6jv/K/xHyzLbSjj6L1vlGLY4yN12n5CS
PeDoEYMEFeKemcny94E7JnvCF4m5Wc0uNdn7p9UNthct+1/tv0p55/vny3Zhfwrc
vnXJ52ilOu8vqgSWpfY2Dy4t+TF93e2OhvIXVlJUmufkYTAIWyfgCubMEmfC/iIN
Yv3tNJTBFI37dlVebg2g23AQ7pvGkVxkr3qao+C8qSwj/J6KvMBxLXhJafsNqIIl
QLuO5Kz9AsUny8Euf6ZqcmAqLzkNJiuH9pSK3DuaAQNrhlylHiIwX3any/ZFojrU
bwIfKhCU3foqz1dVhQ4b1ph6lej6BEZz/P4Pb2BMDm8hN2pGZn5TpkTGd7RM5ZSK
KQwUWFBC74dc0GJTqc7bFDeAudcFb0cADr6jt264F1GzIkiDNQgX6RSf5pvu9YkG
FOTf6znmn880mN7SpT43LCA4A4gMGj52iBW8sdESPPbLnAbZN5xyX7p5/Vg+9hjf
ygOM+vj8zYg1C6awNOxtTFfeV1/CfzS+sfcO1PM4RzDcpJ0ykCJfezSINIXAzbV7
bU/qpkRXfsgxqzZkmO1WBZy1a4Q2x44rtDKKCKr8A20B/39njR0Ya8E6cFP53ulf
c6zEv0XlG6spMNwNUb3KTnSJ4GM5zrIwvmyHvEcY4H5uXr9OjpIttOVu0yFwb4KI
F4ZcYyAEX3KBqj4EeOG4atrZv8B9OD7Va9JHcD2YecqnD+81s0bAwShqRxPvLsBD
nwVu3N3V8RPMGIbY/QUiHxDULD/KJUy/ldRb+c/vOWNUE6t2i6Lkcnk/tgfPUxMj
ROx3nNtCJSl6bns8ejEWBFZhw6wDNJ5W5UjwVGuMR8yKZENNq1CyJ0MNokYUQ1Vf
u5P837A8aCPgW6jyr8hrfqWQitksQ+8FB+7YJTGkC1NSmmt7vZlRy6I7I1cfSjA3
Nguu19d+yNTCfP7OMQgce6NuzonMxPJsSDgZgw6PwgXWO78g6T/vqxHWShHXCLYH
TeH0CA0TqS7HH4bgU9ualLPwa/+awmjPh4lMzg9g7cFNA5ALLPWMJx4L6OB9pEJ4
sdpgzSuxkG+6U0Wluq1o+CJOQvCJ0Onq4M1lZM5qlwhk3zxluTU9OCf1/nr/ASyi
F0gpp2XqEuadrxzKAY6yTqkVrkAZe2/jdVAWF2N6X7uYQfs0OFgWWIXK2nUqQFZE
873R11dcXOpA7cqb9eEXrdDaAvdKKTZ+Zv8ei5z3KecgSoFVvMu3CUphee4qknpk
0uyjYcVQK8t/7RIJOXxIKvXr9O1kde9waZvrjTLcsWGamxUGr/xCxSz9tRpvN+ko
Z1kS5meypiLsf+6gCgv94/k/PEoQJraT72XoIUEataZoG/4n4CNCwK3t4uqbstUD
bfBNOxuTsCpPAHUC7EmN7Jp6nqOUPPYwnpPxjjlzA3MSwA97kLP0p0OTItIj/ZTx
9Ge/vIA0mVj2IzdIPLXNt8Rs7WSYvi9NyWb6XdOeUIz47rHp+26dVYqXvYrVxRoR
qAYvGwslDbQsSgQPlNmEIXphmnyyx61TvL82DLfmT4ZZSCaXgBCBszNhC2TUeXBX
DBOrAXiItbBELPr+D4PVtFiJIQQEydc68A6M/DrCSS0TeSb1MD+RcS4nF1yl5VT0
tTNBiiBFpWywdDm/EElZNA8P0YnderMCEQ90kEeaCbrn3wSwxgXrhLs/xKxAsh9L
XR0mBv+3cMnUmcQgwc3kgU5Ayb48V1OpaWIrkKfLm/31SpWqeniotUJMyvUzHwz0
BOUXAamOqBeTPUqkylXAA637tTExcvy4VmvPvjSHUCvsW776sxnr+o1RQlQplJPW
fvVYCIwbC+cddCzd1n74mu00VGsR9CXDKBRIPSDsjOZK7DG1PsJtGfJxw+UHnUnp
56hWQf4GycUEJ7tW5gn6oNASiwtSL3Kgx6PCcwko6sK36Ghqv3PRG1q6/WpCpaaw
m2XTwPdJR2BzleMhkSvx3+hwNnSBsBAmvRBFNDmp7SJ2HYfQZ3fECDMI8x0SL+Zj
4UGmxvqHoFIg3EnsGpwDIFMUArQZrmYx6uesaPShvTisiOKwDJd7tvKiH4MS9N6I
cy7hlHcb0Hh8GzjYwtfTg3bw1xuvbtTpdIOj2uWO0ID99Mk+a3GLC2dvWBIOH/XQ
AFbfYo9DyWnXJl7vla5ae5eHtkEJqK1uP5KZC0PZtIvOywu/UImdnjGPDEqBpWNt
nr70smPIJjITWdzmXdsSTb2x0Cm/rkHGqTO+Hjil8FF3I4kSNeQChRHFbaVK234Y
ZOnX+Y8ZEEzNT/d+mujphCDRzlQJauC7RW5JxOYpF7A5oOr0qCaipRKOyHZaqtrD
i2g6+3PWmyuVJW2om1U+v/opwQihG8xzxYoRMfZk7vdBzKo924Wv2edhOWUCZqzT
6JNAnoX660XGx//QTr3aO+AleXqwxw2IBxoCosVYX58NWhf10VWQ8ggr64qahhE8
CxMvZRkZNCYaRQEuoc8lLkuNyGT5a1YZTidfU6OeypmuHuzywkLkDqn8JM2daF6g
8NN6WtHbd32jDa0LDu++dqPmh6vx0yXY76pXYEdXs12MHfkG66GpJ6eNfeRE/nru
Q4bT4Fc8bYmuC/MPkOBGj26caFxpyAoOMBf/Z/a+mjblzgVDhD1V3gTffZODQrNY
KHKtXs0ijh9H4T/0RGVMyYUFrAaOHhVwctIEyAV0Ysdo6c5LYo021xqFde1nmNdJ
DOunSoABP/rAqxWiY/pP7G0YmzZLcfGjBWoMAIq2aPkX+cEo1iS+jWyO9dvJA4yl
6uGjLN86cm0QER9lL6cxrOsqmU/aqJKfpTsxqRf7GTwHGT9GwvtzekRfOHI7agmF
dp31nzhPeUoMb59ZdpNnxk1c53z3jJsyXHtIXaTAe7/zEX7Mv2s+HV/zPtFvkrJb
YuiOCt4i7zwmPEthlbyaiE+FkkPeX8dMrLPjMyPKxjaP/E3prqMrxB88sAoANriO
b3/V8zAZYwUm3gazv4E5Z0VraUuhoeC3ev+X0dO8Cev1VLIcq1xyMSmDFRk2Uyup
kebTVcMv0K10b2y9FrRRlXdBSRmDUTJC7w/+F/LZWtERAnxJie2PJoMse0UcEtJ0
k8ddqhbc3QFDSwG08kLzpZl9zxzGnFzSDSViIsV2KfJ2nlP6Jw+rTqizlfr7iWIE
+pnkUQtBjVGzu2LPjv3OHfY4Pns92j5iplQQLtSMuce4yPxc1eoRORtzJIwInhxT
dEMC41jqLAFFVffhtRV0p+O+/pjYoUX2yg0hwV3n7E7sJtuZzBTf2/AyTOzG/rRU
c7R+5rN53bf407uP+MaBg7UlFqoG0eB31Qk+A2V8sJnYaSSthlFs/EdLvgg22rq8
VHVLBIk9Ql+4CqK/9Hbwa2wUvIGFtUM07G5uYPmrps2oRWYvVzCxojmF72JaLuoz
62KHsOtB53hXGjHDdkR/WxB8JUfTwegmiGxwLmvkr1nMXnaEG5Bdgd9NyL2pkJxQ
tc8Z68iHVNBLvyR0y9UBzVbg7yqiGIKUyeV3GwGEW94VYgYZR+MCLE3Hbjok/eeY
pQp45BPhEtJeIHaTv8h6q+7SDFR5WX13LJkU6U3BEZd+kDJn0JAViwrJnHvOg+8z
MtZSUL63Klztr/z1jn1JJ2+ojAxs0fxBDVYIEzR5RxyyVYrO/hfIIr1Leh/A5FZi
RGTe0Rph/4PBIBpOZ8PAm19+PF9Q4/MZsYHLY3tW6U2VfHgbFkIY5/xd6qp9Y2/f
DT96Yg42ttVMh029ISZ7xvXZ32ELmhAN+3MGvg7gg/g/xI820CfXFOTbFfOdAOFc
DRNfRfQZfWT/xLlT5kQXBY1g3HAOMrqS12CWYy/p2ZOzMUDsMDXEmdGpoieC1NRB
2fKN8f/yeBqLDP+SziN/VPh4rM0p3DS3ZCt+qAxi8eYnzyg5zJ2Nv1LcDYysWq1m
TrZNQVHI6N5+qbU8qh84UtBZS7bV5zshDWCEZmdZpF3R9FJ9kN/kTG9qa5oNpoav
ufLlC6M60w9xjkpnE8w7Vw027kL4KkeHfj3FsRvB/TaeEjTB20B067DKrq0/ko/p
AjD+r2Evqh/khLPPP0noCOfO2TF8nweQAIjQb3iMX3k9uvpwg1rJYGIMNb8eH1Aa
AHy4oCcL69OWT2Y/vhdXIxFgN7XEOeBHjlBLxNZQ3Xn2d5654JLk/Drt+up6Awuj
TlYF1ZQOQ3awSulhRJR4si5uiuy1QB82vpShFtc4tCeVzbSgfmwdJC9xui2CqeDx
qBWIL0MD6SkiLW+GLCMNAMRPqwHu5GCaSchj5gDMg7NcvxFePnBw6/lSsSEC9nlR
nGBgFRpbfM96BxdSDYHB+miMFMGH+k0MO+ydGJNJ/BvttKf9daG4wgbjMPJmyB7t
9p0SwH3nespB24DRY2CwbZb48ETIySPVd95JKsUq3LNIG/hD2nTHms+WaLQwXblR
seI3u0WpDiEuxIFEyoQu51VpKSlJDOMWg6cev0m0CdiNQO8CS1b5Pup4ZkO1sgWN
8+YTktKac/b4kro6udKwoDxGPcSg865ecDNPp0dq62JoPqKmzmMPLfKGm2qcQax0
yrNYE4fNPFZfXIfIqn8iUScWFP74XpHWAaY5zF2csU86JTYgIKDbc+/VYTXzjES1
95bGml78DIuIlXsf+gIl4agupmK3ZZ3BedcO9bpXBuE78gVpUr9cSoSY+GDmyJ5t
Hw7Y+ZMdPTjitZGkpq/su/LKbnJX6WcAErbo16eqpX5snlMsQnhOEmB40lLmGaqS
T8vvX1mJFGM9Tx6Ra65t4RH8XbuhW0iwFlly9hWI0gEgiP+jUgJhk/IIrhao4iZ+
z8QgqmVB819Y5ld11UZhXLy91xJjlxJGhO1FjWrrbBYyV+T8SqQHqK+cDKCCFflI
QHrOuBpoH1LWQ787/6eBXpKiaEboMI+aSdBm9qTuyUDjFGlHwetAf2H6QaZPEPsZ
4sXOCAK3Ixs+fW/BfhXHzVK11MVqynlD/AiBE76SMNOYv7A0U5wk5T1J0fQjFBEy
xU2y4JiTDL2BY9KXE+sdEJJuXPZ53yk6KWT01uzs0M5Jz+lExyAL1v3NcikrALeJ
fkPUhLal7tpc3pH1QtMfklAldiK/OB0x/e8B+Kt3+t4W/GSRWs/DvqYb3ektaOQY
8TTLuh5FCWjhbhRwz2VaCdc0HED8Gzd2CO2l+mXbNVPVDf+6H67ierRz7GUEI1jt
RdSnHIGkeAF51xMvtm+K/tanGl03bwuS2VpZagEI21jJIj4HyOUOwITNrbuJgZnA
FTYjxSpg+J/y29OAAnh+ATOjdPvAU6cJCGnY4mRcLuazM9LT+28879fAURqxW/VS
wvEnS6XUmz4kvbl2RD1LvW3/f2dXvNlgC2877Q5sVfHztFTb2oWmzVp4m6Rf6oo1
8VzbubkekjgtH8+ewWyY7QapqQTv27R6BK39201elWehcvvklJMknQ4TQM8e3OlS
2w2dWE/RsARomDtlo04Ri4Nl/aL14PlKXy5Yizx7g0+bazd/H+cB9U52oG2b3i0c
dt3Ob22ZkDHoKrcJkvSNEYjtMEnOAIa0QCUGTwFIJjt2IZWwpzSDmsYX4dW3a3Np
sEZLZHoIMsEml9VeHyM4awnBtgkugOQqEf15YHiy0PWWvyt+98ZQrIHK4XvnVMtK
CuxxwneQ1pkdqPInb0cqT3x68mb7/n2pb3EZXtA8LdnIbFlJwqZcNBIVbUKN+yRv
mAnAwjPAt1J+4WIvxx+GXzCmXsKoSUSx5WLDwKkuHr8XWn4c6DtVY4uNluCszkiR
IwRc81c0bCfmI0mAj25nwuwGfo6zbO8CVUgFa632GDk294B4PyVuCRvzz73oo40B
8x9tpXStuaCu0UsxPMdtTkQyCpHmY3ekFVspbXsggfkFoNOCVSVBObOYmRpELpVC
QRPG10v55inI0hf89zyy9SoOEiOPIvXrQCXaxGq3+tuexqRSLZ+GngAfuyC+IuDM
h4qV+hgUEU9F2DAkg9QD1LHEbWCbi1LXcBigERvBTice9RujaEnAd8IIl07IEY2C
yG44NtuX3A1+9vIRkwwcUIcfrivhBm+O0MolZ4+EqHJud5GBjePj/grBfsyGD8RE
dqhYzbYaD11D7frlBFxWHEqoAwpWRLuw//Tv7Z5UpvdabmNnhkBWl+gJ+4HKvPtx
ZPdE5b1TXWG1UuHFNNojxn/ig71DLfkj67ZbWp8Vc+N6VntRCXE4nISeGYDUS3xf
11+oNrccS/+LS1tgNV7EgnwSljwIm9CakTGhctkfxOHmqzOTyAS26EPgMXbJIodn
TKPfS2cZmdBNZBvGbiaYZSvI/MtH8fSfHLEX0W06hC1KHfDGSVMXgQDjx4BCMoxk
mJi2lhas0O1aJRaK+ry16Bj8sTdxL6+sgG6U1uY1GjqL4ChiSsYbf9jc/K5TjJjj
SYA0CzgfWtjnxlf/jhdL1/6+g7hUDBsbgu3yiIIQiItyBWsekRkuQQBcxKRM0R09
FLox1fYFslm/7fNwkpvFO0rtt0N167IPi5DQpuY2mYmmUattbS3L/W+tCvjfkM/z
FzcEIe7N6xmv5GaHNA1GoD9OkW9KYEreFVY4UR1qpVnWS08onV1L4fauAFts/bq/
QGl0dDXmqEl0C2pfcxR3CUE/abKJjdI0HZzwvpFHaGkL2UumqDXn/ZXh4a/aqxHC
yr5DJObl2deRqLSqRDwIQdDdUhCFzYnVRMEGvT4+Xk6OC8+W/X2BtzlxksDiamOx
ATMbz3nfxauN65vlf9rZaJdoVDSH7GSPYebPJ321NTpKCGJgSOTWkpmtzeOeiVtI
uNKgvd/t3t5KjSfo17IPg8jMh4vbZkXjeImebrE/j/qUNK85HGsz54UySlBXuFXm
w5obpIqTuvJU82+dUaygiIjvfI1ROUYnV36U3ALAmC6K4wtDF98u1pX+aB4NEddy
5JnEluBIu0/BrrkyaYmRVFInfMs/ADZJK13E2JkjjBENhbMCFnDsXfZQjKkVO3Ok
54y3D/CpDTxCLU+HZewszah2w6ZOHozaGI1WYPxKEix8Vn3eZm8M5DEI7Yv5EsFh
3sl7kU7gD7zDdsLRaTz/IoasDbLNnBmprHVKqY2pB/5Hp9rqBHNhoFrozAoIRqev
+ThjVB2cUGBYI2wc8C+kyxKpDZpd2FVPv4UItEL4nve39AM3qnpiNgIPCDjyfmiS
4fv876S4fXvj38vocKsGzOPky9vvaEj/0eBrDstKNRNLe81aZ1jZIQVTkTygj96Z
jkk3DeCaNI6hqlJu8NdPrhbXcbTpVW+eXk4nybqz3StYbasTf3M9JXfXv+E/+iL3
9icjDjKgKVbWJ6Lioy5EY772z0pTzSzM+slOUYwZMOb+aZxhcSS0sAq78t+gV96s
Gk5hgxXIDkxAID+1gH1CgUysymUY9/OvpGWN6+sjm4p0RF0VZsMOpAnt+7yVErQE
MRmaS1TwEnDqvFAtLmJ3PKGEOMzeDdNAzNhAqUO1vy9S2QBvGiw326EuwZZF72RO
mcE7p44vd9/25oaNfUjMdqKP7JE2U6XMQ9H24bC2z9Jo7v5vx+1HFKzdWXEysu5r
wL4Ru5Zm+cZs8esyEvr7NWCfEt3gRh7VAm47cMLs+uD0OCZOpMWFBotFWB+W8lvX
jxFrIz0u55O40waqUhEGOSChfHGYKEfHPnDain80tChfNoHDRKV+TBnrTEHEy8NM
kkesNOIWCq5bY8t20N2/tcrtv73+Lwf+BSCw2mRkgv3LFv3C9zb+6ABsrQEkZJfR
0PoOMFyW7nlYULa0NapXFzJ7Efdaz0zISlmOwGDfF/cqueVxzmwUqF8dax8m81D+
f7L6/9St5KN1Y0hkF6U9mccjegjK50nDVtybSqczfedqacWPLOHLXJx2yml4F/do
DQZwGDjBO9FksRTxWe5dvC9JH+t0fIA4JhEfvSRKCgv3OWDhZeKgvsDK4oVM0ZOl
hypl3pwGTDm7x69v18mhQ1vgFpznAAT5qCfr6bi3nYTJGeAZ8hOw0DkwgoSYg2A5
iXvNGbqJrnJ8Dv2NfSyW33QURTW3AGM3AWwzbErwv0n5kiNECSHfNnwV3O3vsFcP
wwrQdIWzzMO6yvtfw8YPQ/QH/DX4K/LKc6QrLpn+/QP13eDu8O3lb1TAuPajy32k
EVISO0gZvboWczCRngcdqKAUaWtQHerNCgFCjVFU5YaYeAsg49LpE6vmZf2bO7yC
eR0bWcutrvIOTuhfpxslzPtKYErJ8SvE0ZPLgXviy2jBdsycY2tyvSPMZJzvD4BF
oQ6zBKNALC89mJ29EZrM8Uwy21CO1OzUcOPb+WEsvzdLaOko/6Np+jcfJ+1kmU9L
uPBd0shPfqZqpFvcyGFYvu8U0nxC3cBE1BBvBailk+oIV7tP4XcWaJT+T9ggKCEj
33HKZWZjAbXFJh5JPIIi9Ycn6EOBx0/qnIroyk/R1yCfq9bbF9dWm6d8hkOL43GF
zyBGKuniG0grA7Xv9fZrej3aI/AuxUjTLmg0oapw6re4Aw7PPD7XHQmJ89MNn3oj
woWfSZBDicuZvGOJ49L4EdPWMRc9Dr5g4qaT4LizMSPauEGAIY7lKo4NG9U7Wdnf
6FHyIIyzjL9HmtmT/QAVoN6WsnvUbwsSJrMZVIxIsyKMwFcl47YIbz/6XjHCImvn
JmPM+ejZ3Z5osWY2TcmBtH5EvbmGQfZZQKisDMLhWV7gIWW4WDUtIzEgEcsjtaHn
30LAI85/cpKTIrr+DYKqT6JfPMISkCOZ4qbjGy9gOohTtisIyx7QZFrJje08L1Tf
pjdyHZpualI7Q6CzKaSqVqXA/tF5cDn5l7VvD0u9aGzBSTir3S0NK3i8V0M6Z7g5
02UCy/0+LMmwsrjTxI1wt6eq57w8XLk4jbemNEaKiXkuyC+ETPYqwe7LVG+caWrj
gWOuswWFSk5PQnn8AFCIcMUBvSmriq19FtaZ106fxYH94CtnBpdfAzXe4JlbYSQB
aF+TysmE12qQPQJJzVag8b86WmkdtM/QOXlpWoIQPILERLRRKxhXxDtge3Q/CGP1
IRsscaioOpBEDU4JL8RaGITiCrQh8byFYCzEz23AH1f23mEQBbvw72UnmVSnmrzr
qbnHNkJ3ZmhsQHJAdHAsCnOR/I4khkqMtz6fYjjmRo5GAJf76sCoF6NS5sJAowCf
zQ2dtmna/HBpF91dGDM6XomJ0fw1NfWpa9quSb72kuO/aggLOaybtquSVCNTHDxg
ItuYaNMiL/hdb/WrhMRJPhlhJ53kK1p6T2NiyvL82nipmbdP6mIVlWUHqz9ywLnV
w66a82R/Pfg/Td9+59lf2sC7qWdgsWIDZISCGhZLMKVBTbOU6ObLvrlm1beiEqQP
twvx2+DtRk4S6mtSV/RnV8sfs90o1AD+Ho3T1UgkiEm30efc0DCkMqD9kk5hg7Ls
gCFBc6F56L8tfRBNskPJVAhhkweQX9Db6SsTKgRWzscx6VBDTCNMe4K4dXg5w8+R
cQ/F1S0iUKlNjCxrjuWzWYiqVvwjBw5uRDPdY7e57iYnIOVZPDsplzfBAI7LpCA+
/VI0BqmlN/LdNCemfi+bl8PQXzasJxm73z9fXoqCJM6xG1VfFTYds9v4SBuRlkSc
QXLEdJBfOu6CMe8C+eDC7APQ5X9iIaaZyZJppmS8cltdeSshoLATmZ1K1OmSolj1
TzZSiuhwsCuNgi/tr+p8Vz8cQi2L+dC5dFjAeCEHyjKR6W14FqCiqTy+TFkcZ9Hd
biQ5V3ELFIpJNvfjDEK3dz4d0ZPPg+m3pk3dIM6hy23+Wfc2BMGt8YRo/lNWpQit
EvOBhPZfeGikcil4ujSyscpOaNNVER00f7rCR/0hb6RlJ0seLTkMNGBZ8rzux7Zs
evgsjh+lpiqKzAba8dCSjA2Dt9ZpySlfQwiqfumS7ROpTZcuKr7FV4hEb0LCZ+Ad
S0fGiu+I7k+18vkhtnl/P+iixJXZfmRyGIc9Dkz7v9NKxiNO+l0MfE1ZZwf/jeTH
05goowCjy710Pp8RQ+VizRZgQ5zIq92gpL3+V+sLP5GOAENcNuZpgCQfSIsFHoBl
NEFA0+iAzuglSJZqUMKST9tVOQTuhivfi2fxAAhqk//5/JHWz7IjNvcImwBxt3uw
z4N+4js6QUe9KX0zTR8NwLTUa7HCKBaLNHsHZ6NxOpnw9hz5DnKPfEBRkq2IoXJZ
J0id/pswYMGU8ogSKnWYCmbiTsuKG4tl1rfI5MIQHVfRWTsIRIncc9Vcc8iJNLE2
kL81IOwRYUMhkvBOPQ4tiqMo0urhPpUwkvXvW0OfZfjQNdx0Aef6jBu3QXOdQJGZ
ZF3v+C3C/Yig7JawF/7Z7MxGHmK4f6C9oclHezAujGDxyRC/HXJa74gt2kadkgux
o9H3v+3AER/XHgscJc+d4pmW2RDBveuwSOIqmdRUuMlVC9maQkIymdW0CAiJ2M0h
8TrtmHAnaciUcDWqoK27ggqA60YStGA8EKeoFlisZr7eviUBpSjx3sQY+vfOfv3c
9Jhkd4BWhs/352UfMPsZQnA23nHSabOk0ugb35x+uXwfjh4tA1fy9NArK4OQykfZ
7oGhqVHVyrrzr83pt/4msvGF1UiTbPRPD96+6IR9XXZOw6GIfNnH1eDIHk8PX572
zx6ot8IWGYAI3raKkY0kamNB9TgvEQSe+LEfjiOjJ5qFN+CIwzcR/0BARQeuFIam
T8P3E5ZahxB6s5tEbAoGq9/ALcmaDvanyl9EUf/9aZPgxDEA1fLGe2lkrohBI/jP
+Rct36elW8FUU/NTuHAqBJaQ6fOO3GyQfQACkJvrN0o+oXnQ6coR5FMD5UUx6zMw
3Xv0Hsptkb1l1o0vvVr+//6Pl6vZwLiOY0JkwT9Iu9MkTraXNoKseGbFigVcamE3
VQIeSbGoE9gjvnZYoIdMj5EFzFBC5GOLtIWhoMbR1085xla4Ggay7Olpj8Ol5eEz
YiKEYIBWO4oRo5M+s13SbD7K9xj0rw8h95ZJ2dMeu44X5SK1gckWItzvQRSt8OGj
Z8CARZrhIiQEYJf86kmxhco036HaAE0Eex1XDpg4zL/P/d+nCQM1EispCnaGkIeX
sR3EjHSH0lze4bU5pDcJvZiJdMd32EbLF4K9wtdLCZdPKcW+7VlkjmocKJccl8V7
fa0YN5UVZqvAlCZkdZtMfReICI0Dagaab2BnnLzNYH0gucWAdqdGQff4ZWiLZD/r
skfPgPB1IOJ62h5UAzvSk8ixVn40OyYwRkDIofoyYVPk+9LlU94VNXBITCVYA3+i
vwYLm/9nzDCD3TmWtEGusuTGR3y7LMui2yGNc5W2GQ4XOAFXq4S9BwoENgVtc1kj
wtFFCawcfghyVPrnH+ZSwoEYRw1TX/qM5TbtEt9DP6GJ1FlyStsJkuIRNoMuZouX
LeaDcYe9X+0NfMDqQ1MjhryiiQkbMp1CSYVSKvq6LHVm/QcgOq4AVg6dAkhQ8q8M
ZdUKDmawyUon/sbnG+FoCqi5oVzOSGCXmiY9B5UT+BfCb3Rnzw8++mySjFTOm36U
A+DkhNqO0/hRtZQ3YDAs7r1lmH9fi+MQdtTI9/LXlt9ZvkJrEUBXbDmKMUuKZTbA
h3TcW5O38pAaF5vgKbibW6jZj2e9c7yVFNt4X4aPG429BqIWXaMnHanFUXU9lQ2g
UeWcC6OD9sFSVJQLFD0lFziKoX2jSbeOKOhNtF+VymrheYqQikAIuM2h+4M8KynC
jkrI6rMAQusEpAxI1JTeunThaLPaaci75HNu4qKFWl4lLSNzUAq+09uO477GL1VK
APRMWz7ZzU2gBWVacAxVS3SnKh/dJ/GoPc4ECL0d/BQ2AcSP9Znzbzj+08qefLhi
JadfHHieop/ObGzf6AagF4BOMN//jZDb4pOvoZgB16kpCUn8U4aTYs1+PDi9lkEA
NGLjZpRj+um1SzDbmn7vxd1kPMXKWxCwA9J7+l7KvtH/33jFimMBUmBwTQOAbbwE
dfd01tpv7pSjnQZzYorAPOMs6kI+IRb+V+vkqIchdS/w0SasjpYKlSldC2FMLHDW
HUnjqBCkvLwG7kLjHZ8tz/f/C+/3L9OBLcSGkdBwRn8I5mzbji/8TNoRWb5ja/Vp
BJBvpFuVEGInbOwxtQ4xv2qzK/9JyC27jzWqYTr7lVMhRawqsBKRcKizQdWpv2EW
5tPwbauttfS8ZgDBUJ0w2ZSFgaWjIbH1hrYjePWHDoTyH9fylC9ekSd7SevjjNy7
/Ue+RiE15WZcNJnxoE2esBVSwc+9GMK0m+vXjUChDNnXBpjGObE5qvCDhIHJaTAZ
MQpWrmADOmgkqXIjk9mRbd+oMSMPoPMz84h+7A0p7fcuOxRXpu/xVVmiYkib97e8
b18NM+ub3bXET/eupQqUspvY6mu0nzVm4HpyGr6QDsZCiSaaPcoL4l2SwWKVBrH8
8u52CCx8aOw6wLS2CyDDuhtolgjL5sfOXgD03/wUYiAkdgQi723VxwK9UlPJIftS
7BvFn5mGG87719eb5jx620lOoKHE7U4DSRcyzjBLPVuM83ugP/GgPJpTfFwbou8M
MAkAhnLTQP6HmtmdJwQwdrK/E3cQnGbK2OzhxSSuXqHBK4egczfZ2bWKqclVkJ5K
4zQegp4+LUvHEp8zsTdFDBpuN6Cc9uQSSAGufJtpGnLBo33OwgGge+o3/VPfh9rh
4JWNRNNbOUPqEaBJB4/5LMhHKHh9TW92KNmdsZKbaN3GTPYTZlPajVroKY9Z+oxx
QHCqMZLUu0lpLPqWupvO7Gy5FnbDHlemWCQOr+lDl1tVygZzEri/XT35HOTxNVoe
Y/3PwfSZUHdNOmmX0g5EYMkZ+sjTWkssspEpPDs6GqaNBpSHzhX67fE4tZFcUUBi
mJY5eDGabMqd10/6n0Nw0L79QIbnWlSLadY6UUIFhQYVrxCUlhTjx5pgKaS3NyWM
GV7aVwL5GMkSk3DOOkKPYcJV6DE06SJ3S958YdIYDifc16nSN37L69wjMcpfVUSo
cxXh8vTic/vmGjzD23p2Vx7SlTWtvRW5aZxga9MBAwRDt3uoaN26zG7OZ3NZmGC8
PNaUse/w4mAEs20rR1haIfwNTxm6IDYRbOEKJGzfMQNV2DRPG2+7O8de9pB7k0z/
FqGdP2OrreUxLxRbtreN7b4+E/cDjgc2EzPIl7m440YT+c9X0rFsiUgOo62gBqWZ
IGR8sXxp6/yEPeye5hSe0gV3ZFHP3hb++RjIxWXbooTXCp/rcG9VIJHH4AQPN9ed
xQcwl42Nmy/vaHues8m9bD9Fa96dMN8JyqBPhaRWEwvjExnjXKdX4klHqJ1OA75B
p0wSMxRqbiOOIFi3p95K9lmzjoaP+2xXizEW4Qw+hRe2uzO8uzw2EY5dYTRfYnGe
adQnTSxNPtP4mYFh9yfkKP+m+Yk5KpSJJ/MxKt4kh0sog5+uu0246jij2GVBzXsd
4Jj43KOVWYmNVuDZ2jO+TGBYciGQax/+cBYnN23QzSfe3QhZzqiql9QvI0yH00V2
wAul5SE5lhQSIRARTSEmggA2bt2VQ9/IStpde0tXDnkzsLKUg6K1pDX5D9H9eQWF
SCMAsxQalLeNktfcIoE/PVA3j0st/7xT/qjaxFAJKIcYQpUCHh5nNReN/Ovd8uct
IMTdt8lxOUSDo6fj7Xwns0TPeP8pL6/b0YdhSAPacCKawdvRel7RdCWIURpdI8YP
IdyqCSpLNN0LOj1loDtu/JBWKRUDaXTahHaotqoZXIR5IhKVYako2H7A22ahH2n8
qDzvWStYj/bfdGLzTZR1kCVRacNSGKx73cAPsGDUE5TJlLEHBO1di50yX1xrCFT9
NSfNCDHT0ELZgBUEU51W+Bmp141xknJlmECEIBkY2e2B3xCcBZn5ppDQ7hESf2tw
xr4ePQ4eyDTioqjbuc22Z/dGL3zbgHgMMdyTDzu1HY9+VJAK/nHwI1F7xfSfGWiu
HAB/98nJ8cHw1X/AhFvju2rV//BkVMSbdn8JX8/h4NxjcDrJ8z0qs6t7MwiX45/n
G/5a+fxgub2wsvgDjDJXF/2+0VYdnRNtZnqXKZoY48uy2uuuwAOCqToMnynaD2EK
I3X3iSJU2cD7+5L4K40IQN/Tr/lFpnPFZIOCFx43nmDpA9g8c1qYab/RMF+0D4xw
7EelYpBxd+AbxgVpBXpe5dWvRMaU/jUd0D3FBYqywm/tSI9wuLA7nqt/Zi664Ey5
daridCZW3Vl+Re2A+/iN3WLB/IUlMeztMYYfyQyZ6rM9dhMFI5/64Eoie0huYU+7
jsXCPzelOnqyaGkGpZoNrzSUlL47y12+FwAJVr/eyvpMnwuP1V5k1TczX2jolzsB
dWFkbejKxJbYnEI6q9dmcZiClH7AhZynkw/BMwnr/iRXVBAzO0DdH+03EXozOTF7
jpiSUortf+lBKXhM9dqFSpAiQ4SpghpywW8jZvsSBKV7Dcv4Bx2D8F50Fy2nOobq
+pwQN0vlvCeANlfiZmIeV+RaL0H41+34UWg74oaEjMe34lxdJweTES2ZG4m8AsoC
4m5NkNiT2FtFrA66Xfn/uCKeTIQ5su8htRb9hcq35kCyQWl1aUjuz5vFqmsRNRtM
K3F8pvUIlUxB7/9W1UtWksg8vU/SEeIyt1oAUgFYgTKmxSTml2WrntveNKpSka7y
hMn+xeHootQ95laTcEchvW7qYj3BLmV/crOvHBfeagUSyID69yCbS1UfmjycEPKY
NY4MfavYlr4/PQ+q3orkRcxt5Sb47h0hY2EMNLoKAf1nNKYd6c2k5bOk9Gk2tQuA
746/2X/NJrqz57kSlrxpL8s2Q9KbKbn2uYPEJPANT0NLiQ3UdgnsYAf1nZ0Fru5X
AVIQOuUfCkAxGWiacjt7EiKkDpL9npt1cD2LJtTfGf7083gx5VAya42tjXx7SRbD
KkCR48+HqZDxWm0AQOSNesPlR4e1eTD4CMSIHpptTQcGu3d0PBf2aLZsiGV6Ykto
PsiWJzCIHBBlBmIrby15k+wUf7r4dShSvkgE1xSunv5TKUmI6WU5BmBJ1Zeo4Z8q
iCHM3uNUfL/mkDD52YkzrAkIhpD/m7AM/TpPfy8re8/LXrNqmVLd+3xNYFyF7TGP
xe+Ad4cdp3raoNaOfCChMee8JyOFoxo/bvEKeDVorGei6SwV7lktBI34BmAWIpC0
TjpfWcQ2JpZ1cq1iU5UgiTaZU2V7q0gsOPXKBqjv5F63ZTqMwY5PxJ7zzBUSPqzD
6bt4LbZsBj6162B84hxlm0ekwDCuMcdnzwoBoQW6/6AZ0gDqLHgubbeU0e6w6ndo
l1a3eFabu6IhlPtYDIP46L2E3iSvcB2NWqydJczQzMzRF8G0+45r4h6v38Cd4xHa
kjxR5KbCWZlOfXkA9aLBbiKrGtFchgXNqfNZkfpc6t4SJM1fWAimmaOGI+VuCWUL
O7R/M3B0nYX2Lx2k5J0ymhl7Agwy6H/mS/3eMoYq08Y+1rKJtw/igASWWjJ4mTe4
WVV3wj0HAWjVxruIgko+2k7RKGsdQ8nLThWm+7piFuitZY4eH+k8WQmjVDDLpv3F
1Fu7MKhX0sdUD4byfqiQKnC+MNlNzdVVM7CrNt3S220A5v5rPJZHg/VacszAX2Px
NVfhHZSyb2Z7kCKAiPZIIjMyz6ZDTlsiAnX1T4m7dQlxV68P5TA806u0eVmAGpxn
5WhhNFIIyJ+PP3lapZptSqyDGkE8h7f0Ir/CkDEXcZraqdHbTTan8S+nMtUtjlK6
dWFUeHYDl5UKzZjla65wEs77Ho0gH9X4ov4rVG6aoxWBHXHMpZGq5mIw7Pvcyxmi
5P5SFTLc5lxCI5NJDCmn0edef0WJuucKe7035uM0vLMdkoDfBfGj6wOG/TUtLn3j
9fhQXACTC3bVSsi7x8Oof7Ju/v96SKcF+z4bW8XWtw4kj5C4dYPm0+HeNnaWuQXh
+LzrzW+bmo1YJMVsoxDQnyF1f68aLz0jRGHo52oSQGe3y5qdUd1ik0csuNMUKTo4
AYBQkiQAxVUpDGBO7fo2YTtt6a9uxo/G0HPBta2+wVVBU2kb2Q3gKEIsiCP5agav
LH3VT5iH3Gd1jM9OwqIw9E35hiEEtxoiNZkWsVsQHuEi3acPSfYiazRqDdB/Sp8y
aQQ9z4NwEcyA8bnxb9pFeDahfJ5S9WzIT9kJwNwb8CJjqYcNmBOzwzTI1hZLOxjd
To+4E7jZ2VWaWlmXVmJA28iEOn3L7drTgOeGoX39mdBmBQQwj0Wuu5NZTfBBa5qG
fSQJKm0CtmvdECjKbpA77K/pyIn33KNLJ13ASHBl/ifUC35ajXmuh30qg5TjRX28
frvALLziakHj4Me3HDaTVj1tT7KtvnxIVjUokautrTlPWZY0FFKVaPhBQTWwaS6T
EUlkUImwCPdietK06JI6zrxNSQ2DIN1HJupsL6sNvXRbAEe2m9C1fjs2Sy5RsP/r
KyZsepzxFqqsT7oLK5ybOVwtaZv8qob5h3yxJ1eZjeNQ9FZvHt+KuSCHsk+BVSTS
86xGiEzPgQhNM2SS0veYtdW8T9UfnjR69LjaiCGRC1/yBV/59NIEJo7LE0p//UeZ
xB0/tjqflwMikgmEXFHy7+QY0zWV9fNZAzMlWZVH3RIZGDa449v332UA9KhsN1J6
m/04dXXgnd72CP8ur20+SiYK81eOBZPY+5cJQKHlC6F8Op4f2I4pSN4Fw1GoqEkt
tDlYYw17+4JhCF7C9dQJLK6s7kIDcQZHwkgdOoa+jP34ENfCGENA976/982H/wBz
P8ILay2d7BsyNnKgIBUCLlv/4o2ersMHXM5X4HUR0KM30sglwRPi+mqmHqKoDZmk
5pKKzOemBik5/uZsoEC3LxDTAnPUpU3LwygDMEUm5eH4yL2OiMvP93+dkK7saf73
+zHOYt+I8YJxZpYamDcCyH2XgEAYw7hnVnSkIsSrRZJfHpEKSLumIhLWZgorgyqM
hf2M4AEGmtwWhF2MRzybl9vX/BqVthPgAODQ9B8kprKLCU/fP/k8EGWVnJdVFv9g
BlDgXhVnw7NKt2z6YOXbyVc8pOVMFTLMRNfJGx9AzJc6h3Wk8D10fNKLJpyMQo1P
v44xn3R0uFLfVNqrOh1fo2Qc92HxAopP3GuSLGwdf3oW/H+oDd7u7CM4bllDkRZN
2RXrW4nWZIifidKfAbAhMWmRoRvsrvpJ3ihMqF0qoG3y7OyC6iMbWbURFhMAkels
E1BwpZOGUx3GQqtHrAuEoh/Tsz+bKZZ0SeqtNKg9suSjZUlWTN/r/dhqSMqdumW6
1E3bhfR9ebaDXB8rGf0iow7ChnEdnTKVz+C8IF3TC5tq4ivvNkTPdbZyN+OLaP3m
5PWgdKWFv3lUoSgTjnJi0TbY2b6iukqOErU7rtdqllrBru03vdzrgKzhaJoPEEsM
53DDI5Ubg1F5CEFNsYoc4wfg932p97tU1C+x9pxT+t43ypUBbwn/0SFdG2Rqsdiz
avd9QKUJAlP9Rp6MvLdm85yNDxyCj/g4fyvuVgwH32snjwrB4AbCX5ieoBk/KkBW
UBrwttku5bGNL3mkDwhSggCbkQp3D0Xa7+yTumMVdVeqVDNZ4+mIQP0uydbItLWl
g+S7HccTpZpnlMplDYoKey0rgl4DMzioz3aFf+f2mBRh/ne6Kqc5XC0oLmto2ktP
aAokcItvKaoPY5tjS28byuDWO4PaXrj/5i66ldN+/ndplLz61C+gaJjcwWbO4bJa
/ICLTj7jD1wkA3zSo5w29KGFWnvcOGFqyfMAMvIWU3BlBNEmw3PwGAG5Eb+3ZddP
DsKM/uykTdUGTk+9iqQpQh/ntf8WMu59suY2PPWg1c7c2zGWZYjIu0mhJMrBbqoK
Nf7ekw56wwfVBI4Wga8br8ZwuRdu1z/WknLNH1Nih5KsnE1iOd4nKq/i5uVbj4po
aUvCrHLDZZB/sKA6s06+SbGEKyYniZk7cNGY5WQLTzxku3l20PGcl51eossdlRNp
U7ptXhPFGRtrIbo+zhPFCGcMZ61MCx3DEV+v8I/e7HQ4eVp9dQ4vPN5WZT7AWByn
Sg8j1554OEqjk7ZTbZX+G+K+MZOZVt6GVqn4gie2rTd6I+2R1/uXAvdOd7/NdVEb
Sv/qwn0xVaqpe71tE8CYJ82sD2TVfkB/u1/7esNuRgrSxZ5V87W6zR16RuAfChok
Fnw1iiSeqc5TKNOvDa0PVdiRNpxe1TfL7KqfPIWZFDpFJxwP5zw8Gyp+l4Rd78N8
jBDF9VQ0Mt8kuRg5z7M7tKjREKtUltZFaWKsJjaHHBNaRGm/y6di16dBVRF23ivB
GeS2PeARXjHKTilCkIW7TFGM8dOxqjOn+Ay8YYetQmE1MtUXDDSX6twlBhkb9cEZ
auYc3skXCfYFJfTIVSNmnHCwDwBy74UPfTYxlAAtgI8yTQ2CVqOvKNz1eIBuyfHn
O53H5LUwSqB8eYoM7D9BWwauxIiLPZqUg28b1WefU6xnKJrN6f/lChxIE+jDoI4n
ZxWitm2/IRQha552Dbb6SSRuyIDxEasf/psNhFB15VUXGtZXYWbBnUT76EeeusBX
OLAzzcj7bN40uz0kgNc2D1EUn7Xd3RUuTFT70av/eTCbYmT/x6lLOtrPxlgp8u/n
IS5PlqP4XluyZHJZHQWw4f4jwpZEx9uuG/EtC1zox0oC8gZo0CEEddCdxquTs5FS
BZnGt29IPyxUg/9tCtL63yDdQQtI8h+mwP6KPP3eLLAXwEM58bnadeGyKb7NgoaB
/Wv4h4q9Ofi+tIEGYPi6P4p4R1PxYZ0eiy5qh4oPnuDUzUGcvI3l/p/Zwpl93fwO
HGVgrSJayOIR2Sq39hxGdoPsBEL0XgAFCJUlktAeC29HJIylS146kkoG82Jitlen
H5i4wdmC6Rl+p+kOyjsMMEkeqA7bEfuZYB2ihgBMRdHvMSKQ3rRQWHROv1107mEX
rX/ldBHTLW16Omh8wCV8Gekwla5IMQ5hu34TTzYm2kduLOZ+Z26XB3qwW5qT8uhC
O2MLZKPQEeZdEktrt6NB0ZA6pbr/ARAm2+m8JXzK3BYMxBjwM13urc7eltvz+cN3
BiAYKB0qTV5UIOe0rooVVPWDKEvQHdyLL50ULOHyUys50eJsNH9l3Q1zzFmcF8Du
QD/dQAdAMd3VBtP1cmMCM7f7+Mh3ckEJ5lENPJQxSxVCMw8Kg8jy+jn5glJuSQHX
vfS2t5lrk7MFxwiQAouDHyuPO+2T+6p+CMUTuwm89Qt26AX8pBhYoPkXypGX5Sec
PqT4djNxDey2e6/rAnSMqG7oLBYIkeo4E48QnjQqeyy9GvAZw6MUhBRJHoAnd+a2
l/S8V8vyY9Pi3iMRV9Jhx+24b/TFkeKJvNzm4i3i6qlo/dk4ENdHPMlDKcM53IKJ
qVqqtBHOAYMKYkyObYtrZwdDuoOlF6GLzG5eCwb1YtYPQib99rJW1tSc5UzjpjOt
KcHH4BJXFk1NbCKbs7qIemzGGaSeZ5K1IsexMOWtgRzgNRSeRFQRL+t77a97uAhS
FxfyaSx71ahVgqMsL0l2ktdwFSUS0TY+7PycTxwFvNvb3m0Fkj+OFFAWVdPQBSEi
3yLHR+ftPs/b4LaYSGS43Ul6fEn64aLiATffneb1//FP6I1qVZdDAyWaP6nci2W6
pa1Q/TBIsHrc5K7pxvQkzVlDCtKVT8XLSQsQuOxP5EIiWztuYfw6AuBzjChdoRTr
5W03RzRifijzSfxasuKk0wtg4nv7j0cIGIeYqSBdcasZA+5n93m24S8RHAChyxF7
m6c9YVHW898bpGSw6bE163nsVxyswIt/ytbGApHXwxXPOdNp3nMrNS//761uFa4c
0ZsaQAvTLe+g3qvSbPn9ZtdZKyjYkZVBHWDP00m+gXr8Jhhb//L9zuGqgfIPsAJF
4aMgFDzkcE9N+C5V/UmCCE9CJKqEusP7xp3q9MwHgf8KEq3WNwcxRrz1vvcfLDaS
gQlEDx/3X5l6aMWM8zxkFI2Oxv200B9DfZ/OdLAAW2fns+yn3po206XcYr3YL1F8
fCcKVQeENsOFf0pyut3IlM6SZKzlX4zduLBWBlOKxA1Nd2QNwV97SpUrnFunFDmz
r9q0a6Bg7MSRZtLE7NR17QfSrNWW9Exzc3Es2o7gDIuZxDC+wzX7FneT0+J/Kave
5CN/46JVdUGVD3dgYwDU3sgveC6nFtXTzBL5sBX5OlG6jJJobvQzEQSJG8E7xnOB
468OJwb+DKIrxOQ9nHde9EPSURcfbbsTFwtMliYnKm939lJev4angMezLrJemUW1
NjKHQoyOtJlJwotqsby/SPW2g1xsmmoyPDo4HFG6J+qNwoedtOZChPFdZ5lJeRR5
B6460Gwds0UpfGHHtAhrCV2YaQ3zPLpI3IEc9lR4OiuvQJnfM35rU13xL/IyaGdx
tXhS7/QCgqmbBaI2LpyJY1abgsVhimCf101E8xSMc7u084kAGcfRxF8TMWq8Mjbx
nOZdHaYpYOd8WqYgHL8WOVKLi99GmE6Z7v1Xpb9ujK+SdQThqj+hLIsJguu3qsLC
Tyupijf95fvFdcDmOgvAb1GAgfquQG2eL9VOwfTyAGMLuHCUK24PFatCiin+X4ZN
cJw5mbFcq26blMGF83dIUaaUFxWfIFk4Ih7zJXCOIOpt80YLN1HTB7kiwgvuZtGb
0yMfkjtcJUrdaN2kwCo1H36syv3hx9qNh8FfbS60e0F5kBumHns38tcryNZVlkmR
ZWEk1/lAdN67wNv1qDEZYsXfcryFwieIs40vQIyfQqn1SKqSEog501bWEgub6Wdg
mEfPolirPkR+ucM/qoSv9BZM7gkVU0vkci6JEVqA3JBgbWQSb1NZt5oI95cwwWoS
Ch+KWk6pRpR89vzxnSSm1eUvKyDLZATBwHTfmp/fYfhr1TAYlZpKDLrOP0SOvpFP
uRj4/Z6tceAroFyiGByn+bjBjvq2iMyik04jnmXpJS3XkkGAUQB4nTPfs/neQBHS
gguqy9d6xVZ0p7qgPg4azhhitGks70665z6igfGB+r5v01+9RrzffrZhW9Ztm+NX
8dyqec28i/NhFYdrtBLAG3mJXaA5JN248NvUtyCXzCnIpdLEd73NubPAa9t493XY
6xQTcCduQaBF8EHjEVFlSZxPhbDBrvtQRqkayBrSHBrzXVFORrtWUk8pgnnClNwB
21L4y+ENOcldWYm7KKnH+eDsQ0pBS8tuvX7GYM9mD0Cct2d+ylAWG84b9HRPJf4F
Xi3sXb6+HA7vtxmL7DehtZi2y3x0x8iZEREB3ri6w90bySDmU6ZR++HmlLGhdtxG
UOxUbV+lAFKnRTwdwCh9W2WdHBEp49H4KugqHtdrNGPJIJHKEQTKNRdrSD/f5v/s
rtNVuoDIWLWWlOsXkL0MAdLLh9IdwD6UxKIN4MMbhdk32UVHkPKKY2UvLNkOFGLC
005Eo2LcLWrf2gEfgPG3thowoehlrFLpgpIxprXYijjJanp+mYyNmyzxrCo0oBKl
Kw80TMK6aQqsC7AdCPwIgbWg9ZHQj6OCvI67rWFhDzwzUocloFfgC20FLaDDJMN0
2zMpEIiv8oYI1jOyLwOG5FJigNM50eoD8iFveeBQFUmf40MGR1jIdT30b+QSFtpA
FsbkEXaKw7FPkP24AkZUUmROxpdneIexbGoBikjrXNpNNsdANzMWWIyyHCeFtC1q
IFoyT4xjEzZclSLUebp1cwWBNLixNnkJH90PZC1LIC/Z8bsOwg4hoX3fhg56XwvI
F+XZbYL08/WviGgy/+uMgyuUFS9Jxjlv1qXVjXrPHnfIV9Wj+drPYc8jvFtgpvVx
EUuQff3/eRKzlmKAfB51303MxTUR8dLFVRJ/AUNt8jNqnRJKdkJnaL5D+3EDmjN/
c02mDtzKzkx5t1A1CRJWokoKTtgXl7pmlb10Cn82WCeyjNtasJCa09ipcuof4d09
HZQ9EWSUU1kbQ4hMuPLziVOE72O/zcMyyTeuoP2+GpjU041CeFrWsNg+3hPDXD9q
tSV8h84DbBZMTtuaZ/p62WD71pH8p3bEhyfDRDaThZnH0AlbhCaV/5JSGm+wB9Ys
c8MrfE/8lek4+nMsfdISBRlX5Z0WMLmbHTegX+DNjoGu49dfnllvFFS8G+l6XSoQ
W6g98dUEJB/mzHDaSk7N/iOnfNiCp8ysIf7GMwu7H0WGZC9RhZSoTjMj++BpaJV8
+rrPTmYvwUpye20gduMvDuC14mRPACAhzXDdH8gRYUadJkvVe4O+HFx6QaBSjDcT
5F/M/zLFw3MoplmsXn966VWWkZ4f1e9AFBTmo9+J4oT4ADhNyeeUpmS8liU32Tns
Zz3Gfii74Qs66OwNHBmYYBEcd+YiKHrV9mR6+OY/wg3RTQ0+OoGWLOUSccn9xS2x
DOcrXhcT/+7gb0jw5Wwt9gEsSyFOJdtXbDQQ7iYKDG2ELS1TLcYE7t3slxivdlrN
93PvFJWqCf4yDnaJGQjmnDkSvOw/TqCGmXbxCbfXYdoXDWO3cBMT+nZ9WVkuizPZ
ImlbwyBZ29N/669dTNPWLH7wInEJN4T8bnQH6XYvkS5gP5WCx9eHttrEh8sUsfzS
ZiFfWa3LLx3uzLCY65O+G8P6NqDsl7HjYYWY59f12TEJErnHVQdu1w/NWppzR0td
QL/pAl1JyxAaXvdFxiCN/QeV9aFIWd0iZJQMfIhR9hcl+ySBfqF1fQm94H3pY8+H
G3G1rMb3Tjbp9ol9NughkmxNpPHKZqz7bVHp3U46rKAf2x6fXNXDmi8zrCxAainU
BV0rS55M7Smyn900i8YR5PnQxF3nEFLg2h90WPqRzZIOybOX5Ff3EFbNgQXP7zkA
kUvo1YwMQp6+Nk17P4EMWzsrPrAaN/hAT9ELI97LHbB26w8z6rfoh+WKhmd/8lF2
dcN9gbIAZKod2mJKuzw/xoLwb+jqayROFLk02HgtKvmj8FAff/VT4/zfNX9RebtB
1Aex2OQ4zfDOlb6IfNwZD4BjUlgtt8oq1z+KAtkJ11t60odInyZa4jB6vXEbGjud
1m9xBRsXDF6jC+NajV2b70cUmb7vyrB4Q8moFBPQ1CRqTsUISPIEozu5C+g9uOgZ
jOii+N1LdcqhJxfNE6JslX1hMiyF1XeLDZrm8CIUrAyHyMA/CH0A8UynU0kAkEIZ
O6GRH2+IEYZqwl03KVDYUBItvyhS8duhZ7Q0TWkJqD+DQyoav8kjp3k+or6W4TkX
9UUamzcwG+mkTWyu/bDqOGi0PY3NU9/8fUxwdrcvffG181AwfY+M+2uP3mpd5dzZ
0ZLTXTZUJBzWtOYFjZwUhxbGcRfe28ue6ukRrpnsbZiRb+vm/t4PXyvbKrbYDhUz
zBlLr1N3RY2cIL2icgbraQ57tw2MGSpcH/fmW08SNhTboBDeoWuYwJFKSjonj2iK
Hj9RgVDsUbSlDIEWV9yk6gQjdkM097Pk/KPsbb+E/gcyIApUOKBG6VeccnAHsTX4
SH1kJ/3tQYiAtHYJnygAzW8J1kpBCKsMOjBY4ZGrfkwJ9og1CDpaJStki9VAJ3hS
BA0Sehy5q9xTX0lX0NDLZRSxClLrZEQmHZ5vYTXODE4za5m+Y9bACnkelALNwTEx
Y1Zoh8k8Mg7E83CJvxofscgnrf3iuk7xWAMyU1EV6JU9CSm4FjAqyGpinix/YOx9
UcUzWsI72DIMOGjfwb3SnfXnoPtALnHrYZU2gL+XibkuHTkp3fxIdaSDlLsR4VAj
MGSplkwxH+suM4hvM1Xt4p/i9vns/T6BZkGSv74YPBTk8IAFTPYTljirCphm0oP4
RoULuH3PF5f5bciPUR6iHpvRDO3nU4iA3xGSRXPDUerbBS3DoZ8AIb5HYE0W8J/G
XqCP0gWDFuaOW6jpmGi3kXWhTFoBDvJSqHthfeg+WMlLINS731hw7rs+Im64xDPw
r/CH5cFZ5srMzcw+jXYiDJYDMvB1mZWQ5dceia6N/LdMDd7sHMQyF4h43Zng06vG
rvENy2rtgftafigLTSnwFtXnhTsydTPdDyyjvRKicBlskByNmNmd+i8e+DneNfQo
ijAxG4hOONC16Sg7J7MvYabbErMVJP7/peBhXhKdwLpZ3PVhQwkCjyHogLwLEvfJ
PV4xxh/3nbU2wkTNechOAtdPYjew/XuvSJXlNm+8Hk041av6vkWekk9KCOEw3z1r
C5AwJwYe98Um8SAERs99bGoIOaHzzzKRflnJeBOg9Ni3N4pi211gQpmi2340a/WB
W93Ip0BXFRG9rG0rczry/pT4j4etiN4iMrFj6VsxZ7NRKpNkzGqFZos/DZH8TnDm
6ZXRU1jYcIjafNx0uX56YoFOGKQOcaZfMMGuSwKwAcEg0KuWT11b8gX98w/BCpgv
swZCcoa/Z5fgdvcdK1hHOOIl8tYuezNYNiPQkzZbxKmf84wA19aEEDr4Jy+77j9/
h1AurEsDnelPYHl+S+EpIrZBcPE9vKvDn2TjxtJggCVnz64fo9+/K+tNse16NvL1
OJdTaqr7M0k70I7WiJ58MXXap9Z4Vb6xMQwZ2v2QOaceXlLzOpCbeOQvI3N5xMt1
y43UyhoMG2x0YAmCdDsq5e5nLcHUX8bx9FbNhRjXdJpOKI9Y0HOqxuWtUJVxa+Am
Y8z4Gx5bqC5vqgYb8pdPogxk7e4A/DZTDLQL6e5j6uWrEDMu1+VaHi6Moldsnv5s
xOcX1Eiy933cVCEcwWlZC6AJY78qey7DBeqCvHvgDoyq227k95Cq15I2ru7qzwtB
2eP9Ay2kv8S8mv0+rpQRz2jpXm9bVhZqoOm4/dSaO1tw6SgYVK3clJOpPJFUvupQ
2xORQv+T4C6Sj7IDe+tRqlIAiQyPCvcJz944jw1CPCEnbqNcVh/t7ZCQouC9yl+J
es1NVnB5wfCFc5kJogJkGfhfKYMSYPgFbfVUhoutHy0OQzNBTYHb2P2yaOtiYg8i
muIuzdviDXK6HwFmPhwdzcMqaZoS5do5cf77duz+d+FSrgqW43oleGzBn6P54ipC
T3ZQcgDt+Z90CqspN3ej3Z1fxfd6oAscuFqmZUen18r62cgtFI0kCNoDWQUa8KKz
+kK6y/B4wJCW6rtxpmc+i4Ze3DFY3ZkXhcNnpfAS9miL1S14xIXkZGAyOFtoaf6q
FFnnG8ZVF6prigPKFeERZ0rw/mdqf21J/KiFWo0qVsjIQ9ZgHzYYcfV7gsskLTO7
tGG2bGwXF+GN8rTDmeOM+uenLFse+2Kln0AgT5hD30OHUSZ4dts6hrVSFMFUK6gN
wHqRrBx2Blk+kPN/3ZoWzukdqBzaF03IOFTZ1cvRuTSEdLNLUsfKGfsXmOTR5AhG
E4wNYVU+TkYJneb1tjyscyLDliUy85pEDBY2C5EngDY71MPEk97AvFu4VaVc24pk
L+QM6pSVhvmr1NoIszQGViox3uxaiAhHTK/vgGg29xbnM4cbI+LbuQz/GdWWuwUz
9reZal9LCmqF32irEN12PKCqLKI6Y2DRY7SIBLa/86B7Wd1AVxyZ+yqHlKpGWmxR
Dv0qEVDw78so1gu+SALEKS6axe9BuQQQw7n/OeVecWlGPIYTFl7dO/vP9fRSY7cC
Rgq6afRM3/jjL4ilI519MHdI4Ox6JVF/6QPRAhZs2rxdYDnT3eVO2WdfcmZjNOD4
sPT1Zu4ccVYBFwOczjTJSCcEpq4Sm3MgwvSdb8LSEjOQ/sdEVUH/thQRl/E5P0Gt
8h2Lx0fWP8NW9U/Cky88LWVwSOmVdEiFFxGHW8HTo2fL8ypMnIOD9tuPNhtdzFKL
trFzIPIdWMGeCak0+MdmRQ+5lWWs30Q7zjPFRQ0y9L6WsvlOzuNJtXLkI937F8Be
y3hCMK1x3V4nMVR0GdjHZAoWAEABbGEcV8QKsxzOjHqn+JweAy9TxtbGAuE9C1OS
M/YRVs54/2IGd645cnqnNNnQGDdxCy6T7R75uT2zTSYBsE2Vxze0bMZ30HjRZe+S
0VkduOpX41T0+H2Z5jgja77CyC7cjT6xO3WmoIxifwZCEw1qZNrUw0we1yHX6evX
ggizAuZi+dI9ZzFdxfrfVhNr45JRPrKKVRU1VE1XC/Dm3WkuOPgBWmyTtJirRust
ElBJqhdPJ1IngJY+aYmKR0VadjtZ7voU93UWX1tOaPgxQXHExZ/nPp+tvoDXILT1
uyQlgzCcI/5WpgLxn16EDhkrYsNHFJeCitWTPYfFjhR4pkZ1b8pIuX57SJc7DyNL
3c7DktxT5MEI1XofvFohfHFUtdIWgNaVmI0kn0ZZ5nnj/a1kIwFElZMw25ej3HH+
4TwH0FTFSiRci0GMbSK5WDIO167D/Kj4xUU5eBNTt0cqYtD1JpfKwA7jr/2ksnUu
ktrKIIEqCSrlsewWoRofC7X/DYx5m2mKsAVg/cxciWW7LWSQcORKMuhnWdk4J/mn
be67heooEGbx/oefQGZz8MhXbfA0v7ooGGfsgAqLc15KVcE83hRXpV/We1WT/hiB
RMoHkaNisI7sBDbUU+zWNac9ot/nV+IcXXyoErSFh1ZveaRUxCVuYSbMffNf1BbM
rLWR81ioW1t02BPpsKhEHggplemPvi7sIAuZDKHDaBOsDU1XAmeTxiBnOhv0GRfs
xKaT4Rqj6CUffCa9Wr8GdwEw86jo/UDLG780w4+hAkO1jYNEZ1gIHX4AgbDUUyO8
I2rPpzDJfe5XfaVlKEUHBazKJ0vsQdav+3kDMOHLWAz6QkGtjtXyv7MF6NPDIqqx
D4gGSxVTZ9w6VCwfDpXRVUbdprw4oKGDzopAbf7dkG0JT0bx371WW5wCs4xrd75x
FSZgziZ8myBiltJjzjPGA4zAmW4hhO/vyWMWdncJ/IFxaFza36EJVsULgdZXCYKb
pPBRp4ER+zgLuJ3GHbmRBnORCWTB2rr36DauVrsyN8yo0sGfK3VcbNbgSFMqJa5j
Smlt+A1aHGLqT+8snr0y/U5e2y5NGmBXTNuefrU0jYmmiK7DJXlQffdM1Dxaxeqo
QT8A6BjlhETL6F9eSzQF2nPeM2WADMvnsiud+u8mDAp/cjXRBrzWBwqNEZlG47Ur
5AUJwbobsd53LGUAYQL3ATZDqFse496dwTMOt+gQv6jOfVvJ3EkjibUOHz6gu9wU
TtEg++xvq1QxbzO15HjaSDSHuuf0WRHI8QU5juqFusG2zN24NRspMZTSKO+htVNy
bQs1udGbK6ueHkJ3NSBjSuXof2NVhqJN7jkT674gCd6fLOjGRBfhDXncxcMEmNCe
WjE1NqJV52j/abIFuKd8RosX7EvTCq1kyerxbTvHonx0IzTRy89+qoq6Y23g/UDT
LtKb5XCnm/6IpuUIOS2OizLlxeoPA5+ejOwjWEqbDYLQweCONXVOrYgdW4shhObU
GJ5ly5ScYsZATmedDzPJLlY98P5cCmlHwakwji3uRDjgdEdOAjw6CWsOed4EclKe
e3SSH0pA5Tam631S+LkugKgl5dC7tLrnSFWsMOLRv77eY2reGJkS6WGmw9Vn/Ac+
9bEgdoNzY80ms3OukYwk6ee6fYp0A3WtDlSAlTsXPo/93RCPLkP6EotmndY4aAOu
03m6Q8xJNhVrMWDzzyLr9DDlDkHLgP5ea+RivkgLDM34asbKo82uZf6MktUznmKb
3wonaAYq54neiWint91geCeN9LHbwBE1uYIif1oqjXzST+4qr+lZbhdLHnw6p2E5
Zsth90icZfiT0s9ZCzv5jR5nUwKNKgNxQObJVDtaihaKGqGip4BMwQwAohD1NTSb
fOBGKkfN2kMPX9iLip49wwGeNCVB757OVRGVxJvidQKnFKGZ8y8w9aTPUlD8en7m
rFk66F25y8aGmAldJsZJpbYd8q3GXLzrcd16T9j/PiKIf+dYIzEYvnptZNcSJgxm
ijf7sheOLrY97TXze6x1PyVqa7LErsa1O19aN9nc4biq+bF6EjXsZKp5O8O1bKiL
ZSYpoKVo6fPH/bHNXU4+XZLViXeM39cZt93H1Fuf66M2Cp3UcActI7mIdRMCUcm9
UHy7tkcur3d2+eSujK9LJse7y+lt0lsrqq+etw348TJY7POLuQPONIhfhdF+82nC
YsePzMBEHySBOtIa5cFFTwL9xtROxkGZhAUFXlS1NwmEECEsqg0ZdDfzU720M/g6
jFJwwh1ZxEYMvBF4nf+FcB4SmPD+y7JdEdOjq9ox+4Cyzh8aNKOEelpjl3t3nOiY
H3ke8ge5ZAR8ldHug7s9pdvFXS+gOhgyuNFn+0K/6Ljmt90/vRKhPojXKTDszpsb
kAzsx6E5tiuiTl0a2kMgTzDXo1zdiTI2+3rnkV30EVrxGsccQAarcDoFqiz12TVl
zru+QxTa0sBrLP9gtzeX1XXXAumeqsOf/tZy8IWkXG2Z13FNHM0w0QlKdytgNdAS
9cKvzW2Mcv6Dv1Tc0HKvSd+4aWwUq4uRmk9dW9lL41eK1RVO8nz2Cm/nbIBuR1eU
6D95ONuU0dyWO1EmFO2Exm1EzT+WLWMMsTvzOPZA2aK+vlQDAq9GjyO0WyFcWejg
BkaqfaCnaF3EOcVXnmvNzexFBoMzksy7qMEt9LPb+07HrwdpAjeo1J0/u3O0VU9l
MKY4Q2H7cXuT8hpHXuXYOf6qs8svJXWuarve/HVVwXmnBDS0yRKeIXJnbd1pdHau
Ee36KAUmxEA/BZ8kCl9QuAOxCF2VK1DpplX0Y3pvXJBlyJmIwVnW/c6WAE54Qw3X
yLiPCwBfYQ0qeOCesgk3eR2fQtM5BE0d+Mg210KzV0rGhnXTJ7Y2nAv+NWm0f7l0
d2E8T0icQA5Oi1ayJAcNpWxeZH7cK/LFLyqbSbEgEqrfBP4IR+F5IxQfgCD1xFNL
7WVTM2J6Pm0vgHalkR43+B5U+PIAR+6pibmR58VVdxgfNFiEeXlRP7pnfJOoFZgM
7FON/NL5fiqEre3kH5jrJvB+4YrxBmvSRger10uKb+vy2mNoBq7rnkzqT3Ks86bt
12l0BTjgIWaKAT9pqAS6AwOxH3DX880aoXpQ6rSM9PghmgX539t2WAq+ZMs+LEw/
CDZYD4O8vIU1HXKOy5HKYe0P0KXufbOxOKjq3W812qdNzFwRCnBn1QK8WHa37ONI
E34JOP0YyeiEUjnIl7unoWVLFUUt4tRRK41J22KDZbNNIzJ36COb58Zo4UI6Bbiv
EAxczVhghgotN2X7icw4uTtRU9UpciWBCm918OD9geQzPpE4o4CrEM9AVnF40zrW
3GXL1m2Whpi+SrMBR8Fpen0aIuVYum8XlvupDoP9JdiyBc02+INtDkjS7IsyRrpu
BMXx7/LNzIORmAZaK0GwS+s768XSlWs9qQj6P78fTobw7qo36BNtV8whY3GFWoXN
4swl/+TL2GT2bETrC42f9ZDpgCJqyGszgnDVkEKdQAJccmUN1F1Cpth9GXU4InX4
Ka8DG0yncYG/IKZvuIK78TrWH0nxzPSJ+tC8YB3Z1oKNstzPliorblR5YBwksMIC
Wj4+BHwexNM7kMnLvBGAmcyiE8Q1TSrjUb4bG2s7VmNGgME6Dx5cKWK0CKF6fL0R
WzoYwBmXvQoqFoygH/HscUWGK1u/4Ae+g13/3D7vRUI8jwVld9PJr/bupCqGStEX
oLNfRpXeEVhdWgXfyTeVBWyLGWbxQMMd8uAoW2O0nco1vpP8/R0u1M1nyjrHVbBD
lps/mdxxneXaXN9S/DYN6zlxeM9wiKWcuE2p7Vgody0QjgIFYP+Y/wSRskec7QvE
rOkWgL1wCXtrmaOKYMr02FyVlqG8FvTEMUSkF50ZEt+SOQM0Q2D0yjuDbQSJEzRu
8KO3KcbBncb/do6QzAQYMO+4rB52wr1r6MeK6H+JTKFmlP9116MHcMRcZxfJz+4e
sxb0stA7WReqVFaa4u2NVB3PPZcItxXy9eVVYjKv3Oxl1KlBe8KI1KI3125jZLMR
H+Xq0PgW7kTF+LIzdmhLt0Edtm4lsRvL/t4OMXxlHba5XIZEh/9CfAtr1qIC9COq
XNui5X9RhABKqrzrVfmtItpfGqAzUenpKw5nfHM/wuNhEbbizEsCPX6bzI2/Wj8e
xxr/qdk5lKcafwEB0ZXRcyrebYHpLPaUTYI2NRVTfTUS0YPgyNGCFF3fKHir3XWD
yIQayAqpOuFCaQRAb0FTrPux+lLEX9UIaqxMM4sf5GBISHQqbtAUx/+rlN9QicI+
Ixfs0n8cUQN9TL1Y2grX+4TmYfXosnvVIHgMsTg4dcPVWEwAE/KAAPizgQ2GHW6f
oXBZG8lY8/MS5agSUtI+G+OhX+6O560XvxslZmSo6MKdw/XxJWnRSL8d7sg/IzWI
UHra71XY8E129NpLJJm5PTO+V2aM7LLsDyuWVx1/kAC/QNMuKYXwzjqsLHgV+bX7
b5UmpU5BfOSR312okP6KWJ4xKPI9btsyZWiMNaZ+txR1TN5rvdagxZJjerK/iGf+
NJk8BgfoY0ZTU+2DwJWOkbiDSot7r5Q7202gduS9g67uYJ05YhCj3+Xnuw057yqc
RYv0FgWPPP/BPyppWyW8ZycTj3yIPb3WwGlkg+TQI5yqHG/gCZfzG9UAXtMYNQRL
ksJCYvRggCWY9NOd7Vc3W3X0+//wSfF5TNp+vlOP3dpmyj1BZucvLOKuFsCugCXY
C6obKPIbTIrO3T3ECrNZ3wRjqH9XP3ywg1SoGi7zsbgRli2ByOSaY+uo2w/z9YYE
X6QkcdIGbxhE5ks4qL+obV1a31IoRsMPb5q3xFL3dxLZFsnE/OXhvVrXQEmLln/3
26vFg8bT0Ifhc4H2WjGf3j61O5mDi3qkvP92rWTN43W5B1aF0mCiRdNlpTfgIxIL
5SCX81bRXtKnW/plsWuDOiwmq2jo1caw05wAR2N4il2NjZSBYEAEqdwjIupXYk9+
zeM9FSnutVwwATJGpnuexCTACq7nix88N3zI1bWSX7xFNLwX+B93cd9Be5WMh5XJ
HTFAIaRfeI2GzKT6MlDCva+UQOj4vY69lM4304HeJWwAvyVVbduuBlBA48wNspxY
dMkD5MSi/q9QcSmfMfSMPVr9oKXwsj1jqUjV4cGksgPpLWxAlS2FZYij8XKWde7g
U3WFlSJYYV3pEyDX+kT0u0TWi28lQYpbyqYDhF3C4q+q8+871xVxOApmN+nzlqsP
ljT7YgB8XETpbGus10AK9H9kO1hxD5Rasb3j7ilnacb2bqIXvkISD7qUnVUVYDi/
A05GYV5gD+smxEtrW8wf4IPaYx3oSf8BbguLQfRS/x1LZI5TETGCrITu/zzpZeI2
Lz/9dv3iZtdwd4fENwITV261qedL0ErAKF8WY/LImamLQPM+F37r3Oegztk5EP76
XfRrgT4gTIGZgvMH0LQYQG1wepZvlibBW9J2kSDEi8zYae1E2Df0FidhA2ZczR1l
ZC7R9sEP27UCK6lh774LkXrNjUS9c07C9mSS4K9g1eqDWxfL2mwqWSiCc4h3zl+V
V0vRAIKo08zEL2HpbrEera/3YFro2+VnNsEZlCsMNmif6WXjQ/wqrUOAxWTy9EHX
mqiotbehZfiTqqjiJ716yvKcrHnKOzUXcRrF10hHRoJVzhUqVGxnOCCymCWJGZ4r
BGi2g3cmd+doZ3sxwbdrsxZVL4GpCn/ZUbJmvQ0Q95Wm4G+rc2sLbuSKGewxNFs4
d85bnhEsWWlt1RoOH1SXSCrhozRXfXmtekDoBq6QgMb1H7QNXfTs0bKrhKiSN8WB
z25A0/69muzsGDEXMAzUR5IZe7kkDSE7ud8IJYhS6n2+sgD2xNRwfy5L3P8DKfhA
xrb+ecIREAeP/6mUxc5925lA09PXyNFI/TqK8q2BzvzWBrfVuCZ0Rqbm35v0qqcF
EZGBrKuOBSNUlPQX9jdQpxePau26YwhHZzVLd2j1oqreRWv2Zy/MJtnXpxc9dmDn
XSIa67UefhH8Far+C3VZjDHkXmjgkf76hzQQXVA1GM+Vd7S8Z5Ocsn4El6+tNfvO
th1zmaoOELpEaB1e4jX52m7YUMrEqTjCkLMrY6a+MEFjZ0DxdtbxTc1T2ITHujVi
zFZPYd2oVaoV/GBtrNbzV2mI6c3P3jRAcuKhhT1Kdo6UMfFS9Z01HjBTlDitDwDZ
3QGIOGU47U5T25Y9BGVe20PQ2XTMlUnyBORw4iyvvc4Tlp5V1I+KhZyppc3fkxJ/
w1sDcFITEGUMdb2E7k5+oqnjqYS1wsmI+gGR9BOGYU6gZ7ZrRC7nl/viE9Z+ur0e
5zhMtUnCTWykqBsZDfSO3DWxDci7iVs+t5Bq1jLNB5Y5nPl8KEZpDBADOnw4wXH8
CndH9YuQrITWq22CSmfKxuF4PH+BsoIzFfB0hhDee3Lc6UlbFT6FoGcS/p3olXWb
q1ZpH7JsO/h6mxZBBjYZDBX31L9kr7Bd3FSb3kaXOeW2d4GM0oKHU7rTT+RWF+zw
fCLcgXfve8m/ZtenMO7rncv0oLm1pw/ha9Ucd70q1Z8HGaEL2PlzeJF/WZWado2j
dWC7Z8T5CB+cPW2OhsTxGq5OqVW+E4+ovDm0HMtvI0r9L6c1arkU+igIz3GaG2fz
OLWrlhWtEhqzECsuRDO/+yRZf9SynAMlqPO3eZB4DzExsvB+t8lwlHEJ986jy15I
pL/JJZfvlQF0j9vwYsjdVZX9pb4mP5aESCQ/WrZZahDn+mCaxrT8627D2y9ovxbH
1o2Zc4x+ybyqMrSLtOr7CD6nG7gpGurPFfp4af0AgR6/FG1Ww/wTRy31g2p+sJKm
/YSWIlNbU9vx3zJbHTJHbnSFp1/vmffpVwiZApnbn+EeyqIzJs1Smfh0gIyCfRiG
2ledCWgih7FJQrsZIzfL7tBZ27tcYc2ql+hxNJO/YWXFsAKEYlqPi6kFQiWeGcLP
o6L2R7MgC7s0zdtjE5Z8JH1BU9hqCQiP7aGbXvLiYupgx/27ev09S1vdnbOusJXv
rCK2U6/A8C6PvJ8UGHAQ2VaM8YMbP5e9PBHiMmvF7WfC17in2c1o9/oTYn4j/Tph
eVfE92kAKke/iK04rN9HzYhHHOL5fkHtGzRq/j5VTQYdrQrKQRdPmoniF28Lfv3F
X973SVHofGL78mnM+OZztOyUTy8gfUddpbwgq4WdBUrTD444ykokY2eeqRmZUXMk
tNVKgiMrNsaZ9azFYR8Ukwt0kkR9+nyQYq2IhfiYJMB+9j5nRtLvi/dM/cRYDZAK
fNeXXInsInjHXUo/v8NlNhNMtdYqghRE3PuvuSRMhG+X/svz6vBA//2PtK42LPlF
vfP2mW3Yd86x+NdkX3X88fdye1glBVoc10oo0hjBtjo8WJunRcC69QPeYEnObcym
J3Vkmxnj52e/tfCOQ2lj+Rj2IQoUMMVlseQXwCsOfEkhsyzoidTe0EO5CsD99R3I
thItDOome0F9kfLaE7dUN9j1kiluEHIvfVUWKSvdGc7gjddlxskJDoR90Bzm6HN7
J/bwGoHaqR4kzvF3xzj02kmzqVcFlbpJmOTqiiuXjzsfXp84CLSgyPksopb6r0kf
K1ADrhftxmhzbNHhBPN86CX+mu3OAYf9X9EOZkYVqdn9vh9S9/A2aDgPbfT6xoP4
5/OmBomQucx7zMGQ1k7xTArwqwSqJJ2EwwBJ98ClAZTO6JgmAzGZ9VQMSvG7x93a
nuL38pxlBgEUPExqmah9Sn84uK6VwvHCzZA0HpjO+he3nztzt6Nfeum9YgY4MCDm
9IX1Q/t/Luq371yt0fnp8BzRFdELebH2jdaepmuzb9eC0gIv3WNaC0+497ZMRSj1
vnoN0ZXRMstBvfi5cgVjuDz6tOogq6TkwIVP6zWkIHYmexrQnJzagVsFWXJ2Q7MI
UlST1qA4pGr+O2DANTujPrLb+lbJ3H9l2mI0Qs7SKcGG1k2KrjVD3EAQjtSp/v89
YeBS2zhphahbUuorpaG4/v1xAWg2oVH5RFywDC/jQ38qL8Ild2LrWe+ZEJmkzhm4
sygvXZqtPeMnpAZsrry5WmAb5486pbfm7stY9o01t1yD2lEmF45eoCzBjTQ5uMB1
To7wyDrOFkMZLioVfjhQSGfoSULjFjmQQntOxJLa11vjJKE1S+q9z14JJymtuwCB
A+Yn+W3gVedpQyNZrejgUKBjdzCggdDVXsj3CyMK4/g/cAYDxqzJRWS+2JRAVL0F
ibYReGAlJCQNR0wswhYylvRNsod1/g+BEkrS/KRW6qpUE5f9UN2BdoHs5HpxCtDw
zi6Im+cKr2JwY0FwYzvY7f/wcNdouuZd7bJhvuCMYdomfoO8R8dIZXTinW+hB5lp
MhZ0/52P1vcum50kOtGrktZNEZBIq+ObjRzSHPfX0UHa+Z276j5zRHahVmcdzQf7
y2+uuBUv8WhmQhLMELTnpuv4LvtQBHW04NS++mR1UMZsYhmcuokKu9577vF88DRn
upJPxcbZfRwPvdn2GNd79JSNlxL5vchNsPiSgz6j1birG5xauIpYnV9yXQpyYz4x
xmuOFtj6Yd+WmoXEZN8It9jc8trKQCFryhdXVOZGVf0KM2b4lufV+Yj/bnW3gTrp
zs+F0KVzOzaLS6Od2AD4bS6LNAbHK2GE4XHe80Twhpw5EsG+0/ZbYcyGAa7kpcxY
yqK0oIySItLu0u1wbQds/XDp1Zyr4Ryp9TaNqoDBsLlvuLhLxRkOfEaXzrCh+7hQ
gAulhJkVcIJe4kE/mUaEKhp1ul+NH/tIt5zoUILABf+YDz8cykhCIGvpt1XVPhOH
/dtCZ50UI9RdtJQ0RfihSOuLzq12TRwtBb4QsT8ouDIqqlqIAlggCMHZXxnK4zpw
KQDJnjFKLy1IuX5nBJDUMI5eSURojTnIxImJjJVpQLhRpFrk2vTfaJINL5WM3+lr
Kl2KxaEAAetpCIUv0bGoli8uAsEyWo/TFCNSu/W62k1WYeIOT16ZKtPC+f1FT//6
9hoeoqGi5OTjAV/VlB7vF8oM4gpc05798wndJcC8zBj4XypJnkrFbXr7r3WZ12dE
g+H0z45E0j16cu0/kI9zdEYznNNIwwMOCOo3fqP/BQIf8xxpuWGfWla4ugcL/Z9i
Sv8CJPoxDThZ4zJWCi7k7FAnJHD5cLX7nUkolWcuVLmbTwNNLhBnql0h2tsnhTYZ
E4DycjnqwdBBtN5KkIdQzSdt4+OLfwU04YIYdcGXXFJl9N8XJF+V6NdiX59gFNON
vBstKlppqQkfM0TXpQ64+MPcyhXMCDhXdmdb8VW3Or7OEbeIZ9Pm9RS64RzCOEXR
Okigt/GAsEY0BCIo6FMC69YWD0CioF09u8lC1OlveVc2wNjE7maq7io9b87gUAQr
oz/YdEuLTmosMawKwUiJZeueq2RN5qrS2KCT5sJyGIqYlHfswRJnjpkUUDrfZidu
KE9i9TBJHv36WZpG35GmEuryWCzNI7gLrnJshPQm/4mSX93XDSvs1hje/KYt7L+j
LZpISJDDTrsuwXCN87lMrcLYWtb+i3TiJTwJxVeHMGEzBq7FscKDo7o5T3o3aeEo
3jSorWY+l+AXXC+VqRIWBWpa9I8Ue0YtvFRI99bLfVE8vXPhsZEbSB94YwmajQ0R
HPLu3q9ZWzVcMPSEvZNqpytPdBkFBQ7AegbooM2ON7D9DikVv98Cxi6kh7P1Pcpk
YBP1yQpu1381QjwnlM7nDpG1EpaDSj+ziH+K/Bo+LhEef57S1Yo34AIJ0hQUeIyN
s1PQtRjgjVEk8udLEff7f3/pi86hwEtiXatT3+jrWI8WSk6Ucs7sn/DasRfFG9Ty
aliqTCNSf1ZxaCdDlAP8rumFMIi/ygzXfoKSQaLcd+NiBgEdmo5BWcyIwAhYWOBz
VBHUcU2V3/pwiD1ZvLSmPPjiovgom0SUN/LjQhpaLAfyWUv4sX7Y2TxLZi5QC4XF
MT/A3qtqDdKvmwnA0p/c2TkOzSFcKUDink/7yBUUFWRXcMs+olOStpc48KK4RaN3
jl9AfehnekZ4sF57aIMkuUgKj8mIz4VgdvWFV7qBqLmz8002W6tTVTItOljnaXeC
7OJIEZiJNYnIzRw58VRbSJCrmVCm01qAGY0wqmXIx2pIuNNDTBgUftxMQA8gcfoU
IryNU33b4t1pZ194UpH13bEFlKICVbtZ0JXhjT02pfKN3f3LSNziliGDymAtrLiu
ullZuESkiHThhxJ/J7Go6DuNVptPMTR8DVOj2+Udc98QhYAmxTwVtZ2NJHqmYXLG
txsQ0REYG7N1bX4w1WKUxK6qA2TBdNu1WOn9VzJDH4JxNA/zFPEJiY6dHGRMb5Kp
4kWQnTSH7toGjLOsqkxp3DZCYTM41Sfr2cy1B/zQKIzjzJZ0iQeLV0oi8l0CYEOL
xWlWBpRwIwd1rJV0fy0Ss3nthgXZlwjyVGA9EJaSfbizxzF53Nowjrgh1qJwDJjZ
Rvpz/emf4HyK7fLIJ1hSDEMDCCLCGUOvOd1KUK9R/PCgprcXCplloleJaHTxNW6v
y19y/JizxUawj7Z9Vhtzu0QHMtmLjZt6xL6tFLEkX+r8zK9CPdUPTnjmZcTynkfq
jtoFtqhtVz4aUEBdT9urXltFXCv2WhW6lYSZ4NzB+NoBYi+wXfxYArnIIDCDvp5q
7oD3QM17mbDQhyeTXvUVTciLxVyiMdRoN11xiY4SimkWy93RFWd+V/46AMAKHT7b
w18i5GwZgZk7aGTOGfhe8hBE4gMR32IZdWiqC6rbsXB2qIqrRvDiO3q0xuruABHM
laXn9LSm7GtJgGfV2D9Pg6YEtaXewOBIu8sGbtiM7jcHSYjGz15GAOpSdrBQHBf+
c8I0AU7qKQ8UbpN/RInIoub5xl0bOnQGwloM3VDc40bDvnlvkgMhDMlj77c2OnBO
xkZcQqM4GdkW8epMQv0eWX+GgwrsWgjYun+6qmrq6G7pJQM3dS6lmcRybAQx3cI6
zEN12RhUexEAmL3xa/XSLp7b1CDoKJPmvGRjNgNIPJwkKiSLUPLeNLtx0Rc5H7La
WG1gr/kyqO4tAWqa/hsfo+Mfe9sDDPo5syR9nCEAomDA139pXULrXszG4WdLHKud
wFBdbXqG3wlsp7np7RMghOcogjC1Y2HM9eVYXVxmuMVqop7NTaQbcTRKJLO1TJ/h
VEE34ozn4Y2F0bxZpjBWsKktZGhyuD2zcUTbbdosZiQRnWvrT/gEUQLSCpy4S9n4
3fAvpzCHkIdk2tRTCYbf3GOl88P7B0MjJrJKgvOZQ4tm2x/IYlNJdk6EjwS0xw92
a2AbrqP7pB6c1w3dfDyeDa39QkmM72HKXaBgGRrQMYIs0zOzXk5xcNzL7WnGIt6h
0vAoChirVAAEewc46d6mLqwfbFwijuYY0Y6Xy4Wgy+/nxCOGDdoGgkjPb8pF3bQI
qQ1niLlVwLKi6j+m1a6XJDWJnzXE9L9+V+GfieeyRlb6gcRgsYscaCQiAfMuM8eu
NTi+mwvpDjPuQSzzsvLCf2e/SQLozDmQiKQz1ANjazIbp0wZFQs61CUNPjiMfdOs
wanwVgPrUqDM9VvsgGD0+RwD+9e16U6WQ00vs5pz4I2DRDn8bovhWuN2GB5BQzTB
m9LHoCQEaa6HVyDhuF9tYvTsjZ9pJX+0y/7tdbs0DGI9TZN0SkAhNXZ0ISwboIB3
MH9YxW4GxZXGsQwRo0GUJOIC+tiEntT/f+BtmQlCp3iIKmNhm/QfLm8P3gpVjww0
erAi3WNL/hQmqh29ZP1mANrl7FnEOZS3uH1NaJHYaLkphLo8PMAxONdkd/6fqPtU
3ioumi7q6dATBJIz2UMnLUOW3jceLbHM0+M/txXKInZkA2mGPZZqYI4O9GafIp60
irFa3aAkV9mQ111nM+OOqNyoporDAxBJjkDenF8bVKrJ171K/O6FEsTVN4KP9mod
kfYGwkq4KN8na28RvmAfAfinJFCtmnJ9Tm/6qcFoZVQgBqrO0TaywY2cIQZqXQMx
Ab9TPr1gtQpmIHVXM3T47Mau9dd7GTouRDU8cQP5z+Y6g2B/6H7xf+Bu7MFYbXuZ
qYCHKYXBltFQe2ryFn8BH4VOzgsEV8HxdoTporuTH/6PhmwYIPy4+A0mhIkZuO2C
M8xEaNiIBSvlyrUhkxcCu9Lp5y61DwwVLeQdLZ9R/JhnJ2ZelYVQkokt+JCv8g7w
lubuiLgsvJBVUxKvBiv7ucPxAcXThQ1Or/1e8mpQPjDX+1Q0hLa85Ukz+SnfpbWA
`pragma protect end_protected
