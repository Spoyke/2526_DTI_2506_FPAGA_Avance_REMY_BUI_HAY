`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HrvAKrNrSsMyUppP4FIzqUOGlf6+6a2+cYcTWONJPrEV1I7lS088c16IZKu81Z+S
ai71dymwoSY/GMAPKJ21IABw00M6ojHxYqYF5vPxpQiE9iBh9KPj+VVDX3a6mFLi
tD5bqtr7gCt72n/Vh4kUSpEKeAVRsUw+ChwvcEZDt0c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22848)
J7ObD7YdKIJiJxfhtHcNsvXh93bnRteV1WqohI+UCsKZ9oyF47/AxDkrqbdGTupd
XxoDqy6NfGa6B3LWBIEJI654LA4OlJoUM0iL+m59+6PBkpZ6CAn1Kf9mv5GXwNKh
1BNzkdPJjVtAjU63qI95XU/uEBnLuC7s9/TILSCCWDNufcXd4ZcoL0O/ggUOa3B9
5y78SBBCj/3+3el7MulJ1GjZr0nU0bVybAvmC9Re/kpR/4uc/HuW9Oqtp84IvjSq
nyktKkoJA9XinHaQW+ONFdJNMVo7SAEgAvJi9UeXxtIRyjvS9qcQv3FtBhL/TYGm
wyAwJ53TC3QNHuBj2Y5mwSXK/xAhjzWL9sLqM01TgKMjm3i2xyZvbDobpZ55J637
5QIs77x+bC4cbDex1WMIy/VBnBbNK4kzrgUuSJsyRw+qIw/A5aAXZ5Te3UhpZ8Wp
wGtsb4SEuFQTxkcyXJvNM1uiHvlZLQVn3uVNSErn4T6vkUrmhzpaRMp1v17PzYIL
oGM5qJXA83BZSUdLb4Qh4c4ezcorxGwgW7jYQqk0IUzLabMP9Il1jkt7deQTPDqg
x3M8lqN1nCxSwUg/MMQeaT6wofm0Rq2NhSdt7IZRsLyQ+xwSQtlDZyFZL7vLTveJ
3N93uFuO09F1EFSb5WDTGdPqK7pm0mKE8g3r0npb5NYzlyPdif0UMQINi4UMbEM8
sn7PWbQcCxlYzysQ4OC/9SBUaMK7ISmtRqcpwTasL/hltbidncM34lovNV/VX/sG
m2Pwo15/lXO9dT5LBIoLZPyedvmfoBG7noTDb1j9H/vDoWj/6bMMMDSdPH/1BOHK
0/p3i7W/wQ8QGNq1prw+AINy3A5ldfv/v8qrii7kaGpNX+u5bMxfOUBP/kmmooJ6
biLWCdf7R9J2UUlNFPVIRj2v/k/gN0RSO945r1hhAuZnHj04wrS1MlzE/W6DzW7f
0hhoa6/E2bskq6i2YgwDXIjCLX4abvKNpcAky3zgu+XYLWG8Wla30jdV9bNmAfzN
YNC/A6DNGk8MzGnKhQI6h8jIprhBXzZEGTa4drKKt9qQ70JgKjPHCy9jEUmYeSe3
/jiJX90d6AUxsgClZUNxCulqs+P5PP5W7j1RORLKLbEAdenZkXoB8svVVFoKZ3/7
+sozrufKlu0o5gnFLSJjXcBdCHbj8hl2qdXeFAxpljpb+KtBtMLm+SSVib97vQqm
ctnGmDOgwkprynmWOLrubpWerwd0CqXy9yXTSc0IFG2fAMrNdRbOlA9OC7Syw2kj
Kim3kmEnp+WTawPYwdcHZfRILorAIiA1yeROO6io/L6zEJwv8dVSwxsYK7pZLjNf
4kbyupiXeI3hZDk4qL4LDZ7xGh8EAWpbBfm71qUqD5pWInGr6WZ+LMOhhst/aaN0
5PovFF+SSEe/teEf7Vb7oscPbyvv8ITApNO9xUHdGakdaAqOsvHdEs43r0F6wPQ7
y24FlQ1sFVyErplK2m/evXdAW3yGoPcy0HKi233WbPJdaopyNoxB9T9nhni4ALrC
/eGK9SFDq/vrcIwH/hcG33nh75IYOTlz8J6SwvPgDqr6nXNt4YiBfdqqdWxJPM7Q
nAR/xHCbzIX94ZDYRLw6H+LWKaFqdOLQJKd8gwzGesjutdgwk0k+BteXGpE3fFP/
cd1qAGXmFkStmpdeXtP36kXSjTKzHS15LE1jp/zyMrtTaQS6ZshTiD7K+GlT7lzt
Jd6rc06tNyU65eWd5wDjblJzT1d3tqdAMeNQcDbw+glnpetitKklo60gew7KuST9
H5IRnlLQBshrTenZdkRcoEO7HYlDOqdmXfgpniaqM3U75S3JRc9/Z196Z8FjUG0P
Y2Uxu9yzH8hanwSz42N8hnLC9YhSIq9qtvBOC+OraDIaZF9kqNB0dU/WV5ShMqXj
Z/nh+QUSWJQU+IJD6uTgGOfo+Y8BSj5DQgAffYbSxOe+XOHLJyjCLEQ7surdBRUT
k7DPxksvvjJZ24UlZqhpDVhfSyZOiFggmEVO0NeL/X97T7ZRKTWqfcGCGerjERzb
DRHiXIdukpZVXk9dMLTMQPI1jg0wjxOY1/3/NXqkfzunWpQFvBeSjhGAs7+m6I/4
p/zt2eYJKs0c8PbMQUN/wZFVtjgep6vz/qjcSp1tqfzRMFLUtWTG/hd6yj1BcjOu
tervlOtzzUJHRie2tm6xF1TCtusuc/f1W1UlEnzUdfypBHsB7AsG3+uhVySabgnV
Oac17kfiD8eoJLFxoT3MBCPcjMJQXwYdDaPtwfsTD0rJ4O3a4uZCoSmqpVz/HqmB
nk4vdC6RU0KdT8ioqCpcjR+zY/cwfZ4pnIT1B4gZxj9DPYQtpX3BX/yoHllfZW2U
XEudada5eCHmZn5/o5UcTuHxuCv2e3R3c36cjyYUuoPuVFaOdHC10+gTS7rPvn2p
qBJ2r77cnONlNcl+U64pHP21SRmqSghD2J7i7Gep8Bjv3bT76U1MTgtyM8Y0G067
Ukphv84NC+yu2MF5vxqS/TnY9KiY7C9gLjk3P1+d7kUFmAYDTqwLFXF8SGktTY0s
SE9ePK3/NRPq/FEfSAN+/FW8crHykNSiVmMulQw0kVnX1D5uOjOvINAqQkZBGzSE
OqG20+2Dq2V0Pq3x64qqf2oWcDcwIFeP7oTkSfCCL+wIwtRPpFdwcUd+dmQSObK1
svyL5aZqugzvYBUCQueNiPO44LnXJFaRHGLwZxJsfOu7FlhXxbC6T9xCUcp8Uje7
Cua+yF4dg1YmCzgvlYrkDUj63plp201WkeO+3hBDhktebnxmk1lCGScy1pxtf/Iw
DzD2U66hRXzlN5rmyvHt2VLEFDvCuZ/PhKLAitcz1whhSF31eSG9oh10kYZKIhty
icyzh5tB7TTZ3OtCoT90PTFFp2Sy9JKhEfCJC3KilWEee6Z45PvSCbGnOHpsP+z9
WmArY0f42Ycpynd5wNQwu4931IiceIP79CPcmBerzuCUtV2ZZIesxHUbbHAu+63Q
ll8WCkfBNzHuDXiqbAjau4Rn/8i+GKC4K8IB7Ca1FgNuQsQj9/ysm9/EnHQSY5E4
RPjmEjzbufWvEJwEp2CpKHYQcblu3SsjCk4UIz/qy+5N0+ogbjldXtBv5Uzs/Zfz
RUmUvq8XS7Y2TLOazo1pzQrEMbVm4i1fyJdqjQgvBGtl9C1NC+PW8INAPkW99iMe
qUDVdoeAHg5wJjx31TnxrVRUsJ2CUsRAzooTSGNQSWu0R3Q3fe4pfesPgCOQNN8e
EGkP9w7zVI4WYI2X1aTSpxwSl7rRlBtKCBWPJwNXluShCcmtd8s4zxm+wUF9kI8n
4d5iBu06bQar7UG1y7j4WsLOiEYLe9sH3TnJn3/TGtqKfV5Eo567ZMMgaO6RFbKT
NE4ndoy1MLh4GCx5B4EZcbNhjkAVbMLEKCApRDs+NGY7OE1maytXB41ipsWailY3
xMAj4vnhXgCcY9TM/kYoKOorWBb08Hrt0XpQYIl4MMjtwHCB9663dvgdtXlbjh86
OueghI2U10OGYJjoR0uQOOFzGHGuZIeHwlYArrxFvw109kh4nCVoR2rsrRW59aQz
U8qwf18z3LkaOvmLkPcBG4rbxSmPi4CDDXw0zzhK9zwjROGvXM2dXh8XRIB+BmFI
nPFBYFtoYkTcANbricOMvHNOTyw808Zrs6WhOJ7AUAhg2L8DJGkTHcidYbh6jg4G
i5QquYTr3BRL226wafDuczSHzxwoyQ3MZ165kiubC7jGM8kpB876aSrMx6F5mDRq
HnqNqR9xpRKPof8lMYN0y3w21jxxYTRvEsCOriIVA91qTuiXlXL2q8Qk6jjKPGtv
g61teqJ4heWsioc5Re4JjWXBGjfDvjwX6ipHtGfkvawgRa0PvmCu6Zn4sHn+Uv03
iH08v+7SxgU4NCiZTlfAM31gwxf8fmDxmIbZ3V6VF7zuUWQ9H0nSTZqyqp8CXRnm
McwP0oJPfDNknVU5KFdiNmFThw32FEQPH6lUUw4NUxumLHuKDw2CML4Leup5roYh
DZj6DuzoKJNi142OelppMRgxv687q7XQ5dYGRNqZU3fFQSUvz2+D4yGPIeBu+5x+
RVE5g/Kq45gxA3ROe5gx0m2hhMhmXkiX6QGYKOeczHSmAORRah3zVUFF66DS7MNC
sm3TFHpRDcqZtz3aqIwrdASBNPYnE2GZPQL8HORRyHC5bJZ0jQLxOtzbRmBOG3zZ
oOpnSacG/KO309QArdGNBjcDP2PNLA8ZRHfeC5jeiKJzn+O8maRxnDX/Kmi0+gcI
66TF7sUmX+rxYEF0EelOxMRi0s8BJWdLJ1UbgECgFGbCrJEuUMzTaklzu8bndvjT
qL9eSlaaIBNgp9UmkmtJu/Qz3Z0JvgR9Wt4yRU93y0koJtZNgpStb0ACFN1GspiG
abFLoQ3CdsP348iTemHdovnauQTM0cQOvn+wAX3kGimAkgZAfWXsnhfgY1s7NSkl
Cmh6gLUIQot7lpt6thn89EWZGjnUDmpcWDfrxnyqMSA+cbHjLo03zSPg501hbEIE
qY5Z4IVH7v0miaEDJTAAgFKN0xMuDfstDntvIIfxT3vrLlbEhk7+Ua8WZBdke4kV
rwBo2+ght2GMGBxKkOOftzQU5QB3JYwZ2xIfdgAD7w84grDDRtjuN1Pb1t/FniLb
huhJ5r/wzEotZQzcL/TOZAxhdnk2ZH7JPTalwGGWpU4NuTtAx7n5P8F/g7vN/zms
A6jNmvrtmJlQfHix9osj9/rIbQKu6ACAoLH6W+YGlmgjmPQT4MPqpSAsbx05jzoe
jVPdGDoTH1PrvmVsbX7oBWK85o9dlxHTpfD8F8VzDM/eRwdJ8JKSiVr9KWhoZKum
kfPHnehf6j5dWIPBaj37ukgmXydXCzk/MXKZ4GdsqgN0u3LNZ+V91OVufAIiRLg4
YfaGN0I3HnVsg3Q1i98fKWbeNXxYIdIMNF531RmiYkvb07x78TYr0h7qXeUyG+Nw
nVpTDmM0GcrnpjhOS3t1khFG5oaFRugCOD297/RHrFgtklS8fDLTKlPZzhI7WgQT
UfymGJbZo/ExUNRGxCq4zRSxwYd7sPkYqeXgBoOrBXV54Biua7qaM4t7EbpRtHhz
77WXOz4cr/Lw4MMmmp6aCFesL1Hqxm24gwDNAj8SKpKcShpnWTuRFZfbSN8Z2C/e
WNaN6wIcdVTFzE4+Qth3XaLYbJYkmWPRGI52k2EIby6awhZVwPrXMQcPkgtKzGJO
uYZSdyX9HIZPBgEZJljbA4nh9+D7EEiqdy6aAdXjmIATvVY4kWCXrdpW2CJu/1W0
1pmlwDOnDgZ0h2U+CEEdvsa0d2UqRYV/c8uV5QYoa5zhI7oTtSQq8q8fzsoz5xd2
HxM+HzYWQqOsHo7Q3Mr43/QUNJrBFNz46Y92RJuCb+PkAYQFTlHTgCq1o04LuCVK
qMwZ3VJernZXBZJwUV1Myjp2FOWHz9hhyZ7ke0zPZwoKw1lrFpSsIvXLblbjcpv1
G5GogCv0ml/3N4mtIp0qUa3DzEX3VImpEx5cE7NBn5xQpqt7qwi9NqJZVhTAszRU
Enx1hS1VV+6xASDDd3c4zNb793fHc70Chixs5oPWngIDaiZg58g0HrcHEjqH21w6
j5vsFcvoOVNxpy6VMYUpwkXnrpk9gpXbGdz0wMCNaGfOkcQId/nxMgLUY9zx/U5e
H2I9W2zrAIJBR1P4DxVxrFyTQHBBAHEpIrCkt9x7gOV7Cd2VIEgItyKJWcGqz9D0
C8w25l1mePxEVswnmJMhy3z6obccrp1ekI7sP2is/RALvGGNGpUt3GaDQypzzTSS
HaCbsdJrZNmUQcEKrf/mz5Kb61O0PpxT4kvJKoL2YX3UqAOWIbYJeRh2jAMH64Rs
UFJFUxhHgi1lKByWSsp4sv2LJ0dG4AUSgsy9Fih7JLm3yciPdy6KMfv8+ZNr/0qY
sAx7n2/bJJyRLiYI2n4fuzdANtFuSgFMBb7LEpRucSTnVYAZx3HiQkbf+CEof1nW
eFLpfvFnbkcGqiVlbuYoPLS8em+iDyw+/NuHNYJX2Yfyo0/aR/d3Ssi0aER8xP2Z
S5VP4TRJB7CUOCC5eI/TVJ1l4K2uPm9wrbBQOlPZ4hqSX8tpPFqtT03RI32GPmHi
Fv5EGZBomt6/OqdltQ6LsDCXVlOtVFXPW0uTZun8HWxcQxyc3LUKBqPK+loVv07+
t3cTQx6cKP4SbhBEpPG1m8BwemikFm8Akz3WitSW7G3rGRdKKcWvqduL11x6n7bT
ALHfqM3giLsTVJeUCeq9uBFedPbkgoXQ9qKRqm4DaHr5V+4vhi2KxTh/sC3jy81n
kJCr5lhWB+Zt1Dopcy/qf2PU5w0RAfFuT0iTdGz8owN4ETnV4l+398Qdy0SSTcfR
5f2gp2fvi/AdYN+FaHZYOJ67n9G8ZIjQAuXBXAjmglLczDwNL5KtQedew6cfceWc
s7hwMoSm9JuDB7FVXQyeyAnDXoe4Tfxu0Pcg7IVOtxZmTcXf3RvtRQrUSt/+XTfk
i5JBTd0HeEmO6lirbeNr1GNUmInsBICktr/Dvum0ESaFx7+KnJDBxOvrMagnni2b
yc16S40IcsXRTPoMIzO3JtI8AWHbxTo1txBHuyEXtSUAznqJaUNOl6bRDHavDNQj
W2mT4RTuSeSIVVSzlmMWw31hYdep1v87yYDJt/miF+FSftv3Fr9yGA1HAAGXbvTa
4gRutUjXyEkZsJ+qn1c0gguc0XKn2TV8FWcrIdBToo3P/20zCB8agCXImRIBLz+Y
IcM7TRQQDB6SzVRXcgAkltnwqi0gcJHIIXtrwFTZMfvS4H9VbReVBADgXxAWrZFd
RgRGDgVTx1m3gkM0vg2XUF41Nw0EkY4wkigYSRhS/rZPVABj5m93aT8m/Ege+dO1
JU64Y/vDxHyUtR4U8k1nyoOHE4xWJJ2iv5ClYuf984re05PskN9l9hk5dztX9JUx
UQluyZiqKvxoqTUQyMc6tfudaujvpig8efvLluGT24FfhZ4p7Cpm85YluB39Khsj
iZhQVA6VObkBCMkoc5MVpAnqY27d6zwdyn9V9E+Io+Sr2CQQS047AX0V/8z4MYRr
qBt6f/SrmNVQo7Xq47hqk8UQvoszBn3tMSglUB6nX3Nw8bTKeqATpw7vqaXOY7lN
+cxZFl7wnLhARPnGXhsktLiXZv1nWVwgSjisOGecCHHRZQFda/6CTreGSvZgAJXx
8agEeKD29Ww38bX9xlU2WdddmMm0Q6JeOQUQWwAl7A3kJEM1RST5fTQ+AF3kAoIA
1nykPj3vO5IbPUQv55DPBYPHHf+hrLHV2gEQzef6G9xMk5aZMypPjN0z2XLfqtNc
neq5LPSPwvWDfYoExjPEKe+WAgNrAN9VBOiHHr90665D3aojFgbZCR22KLInq6T6
MXe98Vl9bst7ClsbFr47MF6N3CvBip/fpj68BIj0/+eabrZnvYrISWz7yl70bWol
iAePhJCH2k3uKTPxe5ydh2/+UNJF4nDtH5GWV/2X3l5eI0TnGJrdPA8jCVc13G88
CKDLmjBjiK3FoV1bD6AZ2yK7N9auwVCQg1VXyyftlovZaWhfTAGhiDXhQlOD/iV/
WSfP4XVV9EWq1SLC0ZJMJMp3rTqR/Qs/gzKv5yVzTGO4s7MSfrvhbRLSIzDCKB5S
aGb9Tf0bjuj5nyRJsjfOWBGzLjLck3Hs5A/YYpMctjkglEHRMROkDPhKXw959DHc
Hwujb/nCk3GdTD6NhbvxSShKoIepXLXA9UgC+BQdARrqhDfne9Qj+DULkDPSFU9V
07V7svYPKI/UbqiD3+D4SKURg9BwryU6yjxHZrCwLV2nqw5KDyojxbAJtUjlEdjm
sB79V0qeR/HvkbkxFQYM6LSj4FXgIvbbvIZZ91Apo0csTQJaQt+qcMhMAkRApQnH
wzQCZRaPucE/oaX0b5FvAtXHy/jPIeJOoo+dGphqB7vxFTarF2RoMwUDBKrQb6X+
GxqFDEJf1AXT1mUfhJLjic+1r6vcBup/LrEC7hl/aHCQyibtnTHOfE/RxwQhHRl+
Z2zXUYdlDp5NLwwHEdZQaVXALo9ksOk7J22M0A2LtZn2cbo0iR51mcrfY+izBA4B
3lFjQf3nX/km1/F/WAohzMX+VVwxJxtBZUHxw9oL9dxP9nyWkXmUY9a5u9wJM9+O
8eQ5qUDGaqgyLVB89oUIciP2hWT8vVUkIPujwVfPHGbNmnamLwIerf8q0Dx1B1jl
ZY+/g22bH4qMBiUqLl3sQOeX7ycdW8nB41LDrsPkDXYKfdkGkv47ThK/AMUuFdTD
yBa+ZVigF5UYGKhyaIG+i0On4l8yS5dZGw6QZiUnPkG8PRKIHcwJTf2LYH/RR0UQ
nBeWln4u7i3DzUSEn9/OMMbSkJ7qIJYMa7kZh2mZR25dCrhhR7yLVUZkVLWghYYN
H3Dd6yabCp/ISG5iXdWnXwndBVcujpnShgdJXV5Pg7ij1i15MkZa5Z9OX060ap6j
tUyZdIGSS9b2u9+EHr1PtM1MW3/2fXyzWCpWNvhYY0+LHNNwEJSgKdgvVZfM0kQJ
DFzu29yJxabhb/iVISKzAIqeiBsoxflbzFRrUU//CKe9sZkqUxuXOGt6BQkGYtvL
e8ge6GGTvu1o4OHrsySePQ6Vap0DNVX64K55pc6eW8VJc3VJqC5AL8NbhrukHHLL
/kewXEjwyNpybEdAcdI21O15HIhJC2j0w6l2NjNl8ky/WejXxSTHEs17/iQcOyVC
ey/7ukUbpypoAqowyXkpqop6TKLHt2NXf+1oBFwiFKAj1wpW1n7a3xJ4RtW6sJJ3
e7KkFzM4fMVU+rjHtVDjsSfHxY+Cqv00a7CtkiRN4kbzmJRq5+XXK1h88eKn27Wf
sKXCzVMr+cVDcLFxGSs9F6L8svmxnNnvBaQKdylbAZ5xnFL9t8Bq5dDbiCoIRf5j
gBZEpmFYPuCDawHUp7z69l0tpOZf+rlv5FlBwvAWVZc0QyiEAJyX1zN7MtmWRG41
unZ8ZI4d/i8q89bzV9MeserrAeX8WGVr0HCNMyCLeAqT3yb8UY4AHIAnfRjmnNVC
gJ8b7aPh9oST2XEcw/EEUiyx9Y5cFZjkj5rWljLZp41ffnKkRcpeg+2ORs1eH9WG
SlHEwy7g73Z8OYgUJ6J+XrzNgrDLqxFzvUf0wZ4bK+0TFfu7sY6vUmgemPA2T/a/
wUdctAfbX291dLjq/3oWtG0mVdahdDFHhr0KEok8WDIHaxOk4hkgfIjm6hLvss7S
qsitZyKOq8xESWgoJapQrx1uMnSR3a8mSnBJc0qv0/Ne0WfkyS6aa8dbOBxsGhxc
iKkjepxKxqd2oGiYYi2ogBV6oHeHqxhN1yajSkwZYQKGDU6Y4PpjdV8GosZVuOCB
pREG8rGWb9LY37bohW9KxsWO2OoA38KrDQAkr3gjoEqMrNA/MVlacR0pfxJR+k+Z
GxZuKVznXc6pY2OyN2emzofPdfAcOMUlmHYv7iY30LfljCS27jDvT/w1JeQoHhzk
/UrXg+SdqwXFMtyhFn6zNDHtaJiDdVctv4dTCdnK65UYB8SQ8PGW6c4wSlkoS0pd
nlJSxgVI31osWFeG5b5UH+1M38LlOCHKy9mlWzpOmxRe4XoAZuy8uoK6sSjmeSc5
7LFLAy0FhRarcZlO7AtYgkLyzachEJpI7eL2Apom1AC7wBttHd8GiNjGiXmnJkIF
ENqVB8J6r8IFis3xEFiX/ePLJgZDGw6Xmbhd6S4IDp+RmCVIR/uu5AUSO6X+5djg
esKkJCEHMODynqLvLarChPvNf+NxOJXicEuOrobrKFiWFKASQxUJUsP/Y9fkEJM0
hnukdDMEz6yMbUBBkVPoJmCyKtr02dGxj3VqaYYI/13s28pw6RS2HlxGLkh2ks2J
DSBfHwe9WhKXSXGNUQkCuVb5yZ9vlV6SpQDXEjNdI9/ebalkjK+rEdTaRWGfRwVZ
0QMTuwIjW1oUOSThCchiKr0DNXZ7cSkwB1af0OJnKZYkheAY9JqgqKO8DNbc6Z4K
sUh36Ke0nXwSvTJlJaz2ntf9chS53MPAEgSkFT7GeY9LQIPLkl2WI0Q2vI7Y/1NJ
RyxVxwkKoOB2jCoGpmkCdsp3JmoKtGEGNsmtWU03X4930G/JsXCraUiyitltNrzl
EQezpbLeTxtnj7zOE/mEevKuzKd6lKMa3ARRtrFaRtbXEsLp+oJnyBiZ1eq3o82M
2RREAY6l97rjL6qrZ2WYmYZwjZMhKtZb06GQgC9inoGURZmdKM6M+odPhWybCPdN
7KNr1N93vL1rDkyFJtlXwp1AzzxvYK+v3N8pGE8ZgXZZYLyRYR7ObrbhKy0crAkF
AwiFbFsPGQRAtV5ujbY/3dYQe5xwOC+0IIAXnjHbSVfE3V6r3KjsjFohh80lDiQX
xLp20rJyVREY1YUmhqFzun1vMnElwmY5xrikYcy/aFPkhV7uzqcOdvb3uxza5zkX
71N2YXMrNWoEma0vhqOHJ8EEL6oUxut/sjx4TaDq6E5DvPTjEhxQxnGmZ220JBrq
bC+0Xn7ovkR3yhDnmSw1xa6AN1cEPnlJ4Y0PcSuDYnxKe1aBJCwbPyl7Mf2zUHOc
InuF1y2y59Y+CcB8dRraSPcmHqXM2FTCG5OuR6CU9Eqzh2gdWp/OPdF5KLQXAhzk
HSHIKe1rHgyucAreyz1Ij/YxnvzGab3NP8gl9x8O6AC8beBq6R9Y1bBnoYG1BuSD
sRLMP9Ee8huu/0I07k5TCbK8la4Oueibqmwpw0GjQCWHd1bXMZOV3r1gr8aJ91wg
/1Nu1F88B+Mt26LpHp4MMKZ7RuI6o71jSesfXLKe+DuZF75US0d0sg5iSqCYjZHo
Jlh5VZlYpaHI47dTYTIqXQG43tMmZb8MUtjs0QYVPU2OodhQxvfjUgXJaam4wPi6
pctk1SZ0OjpLEW4LvLu9pu9mBWwJLrJLGqLTZcZMM5m8dQZLuGgMeaEydTs0ckPT
vXjTyPcCXJ47uDyi4c2vGUQLtPHsX6TbWkR64eekIblTAnoxtCQKpVD7t4eeo1pi
r8wmmwhqIFJPMg8mcnV/pw5AG4Mrjb/DGRt65EZQXAkCr/QZ4CGVxRtv+z0BZo73
An7U9MQrkeevIgDpFTD8VkKmeyTFrkjr3SxSCba8JgtqX1uUybRx9lajKQXfLT8A
cLER1E1cDojnULnMpFyLUDHwmBHJb/x1J+DZuMqsCp94Nmir1EUtxfjGTQCPjVyQ
RHs9Ju8c/D/YF+fklIJixJRQqBGMVTAkfxGhnLJiDUhReelcsIKThsHssy4v1b5e
ByjzPtCJx+Fkw/n19k/RLONEn2qRYYX5RLatC19A+nLtY6DXlNP2E+bdUxGDnrC3
BZAZy7YVrmA+/oKogLOhkzU6FtUeyCqjhLFvmuPvr8Wz41ATCfen5SlL1KZQYN32
lLHAXnx2nWvEpmhmmGX0FlbrQ1e9ROOFeyvZWLdFwhENMLNEWKoA4USQEY68Uh6T
UiDEhucmHsGrRwmpMKGupHd7kRvyRxNBkWNA5xYhjep+tl/C3vYCY97BS+gRRGqR
PH40t1tJCwTPUuwYMvP8Wx3T28sgk8SjLIeCv/hB9KTia/T4Zsegcm+zXxF9T8ST
4oQ2YnogBY3me195hUx4h92rDjLN2fJg3CmrpJCAUzff34SOuzFlQucxINaA/fhX
IkmLKnwDitPH7JEB01nzcRP94AbMGrjQs7mNMkzbeu/WuuEgfGChYJbgms7kFFoh
hTZ8tvOYV1BPZAS6De29lQDdvL4b29ZYvXapqYz1/5TthwzxHMw00vbHIxKI1QgD
5cnqsSnpy2rAbJT2cdCdap0wLD5hDNTWJpCV34VaM56XrbsqVZrK1lvO9BJI6uv1
uwlZimSsgbWvx03vP1vVh6y/yZxVREznZqMF6WIkQOxZZggmbQcwgV0dgOJEgdQZ
Gyynpf/cmUTGYqHQFdgq2UFSBrCm+m262+lZqK0BkeG3YYIn23HE39FPZJg9Gkft
NdIoqVQ8H+F61HwR7uQ4KJJwPpk8tcSNkUtd3r/RSRl3VROEzIrpNpCZc+PyQgi+
dbUdLughWVLbouMxyVnJICR7BZDqzgOLAVnPtXRW/JNs/MoOf4zgI8WXE0/BTz4x
Z52zvPkd1e7DGAMgJKQtRLpLCNN46mcFLZhRpMwIqZvkew+fWiG+puxmBpSlzeao
cXpSWHNd+/XnWJkIsX0/mu0YFWKl3/wSbs9gFLfOBpZPKEVrjUisNuuWYlu1d4Hr
oe76kbJz/yoI7+e/bbmOPIPiMoZqHQOaxKrTw0T/L+qvzh8fzNjapikXYLpxJi77
6e0A+eOsYd0N4JmwP2x1bkHWXY0UH9EWA6aPhkoqYuRE0snHO072PlX8yFwWUotq
A9y5VGxeF0lVrDnJy1g1y/ifK7AcCV+3UTgckr/1VOZQJ4Ay/wu/0JvSrGOWW9SP
QyneGl2aiQOivgayvHznitAgzprbIHoBGLFK4P1L7wWc5yp1YAib5mvXnkUo3b10
tZnk7NPKBQYsWctvEwFeFGFhGc1tKG0rD6hkimXOZ+EI5cyJbRdFVJcUZOUPZPcb
pSdXzGBg2BdL2gZMvzL/q0fXNxoG2AZOgptj3eoflrI1ECAUf1TtEiu3dMcVKZiD
1a/1mN4znc6cUuj+yWjNyUzHqkVhXyPfy+pyowtWgsy7v6K5l7C2koD04OuF99CY
pHDhYjyy4i4HZn7jK8NaBWyEMUDohZoKx8bcWr4wJXmDbVx7TltZPF5idXECwt15
733Ob4BzrGTV8I+ara7IEOfQh6cqrI8DqfT47OPQs441ngt1gOgQTfbyLtl+/VRX
vbEsfpoaTU7qRMuXL0SqoCvQazyT+scH11kvwdaQghhH1MN1nCSruo0wXOX/wvRB
TJ6459btVlW9sNRZr4liQwPN3IpQDv5Zr059m0QOMzdn90VQ/DA6aa0ZKLiyDzPP
Vtxj24YMJfSq14PLO/5TdS9MvB12Iawyevdg4OtstsHYNRH3Ug79HANugletoQ2r
NTMd074iafaIP7h38JQoRHeILDsqoP8vXwLC0Op8yVYRjtGEUb+TJ04Ak7tXmVla
7ElM0y2ZPIr2ZhiCEXlYCDrTtKW8mP2r1PL9upZ9iccvURJfBgBl1IHti9oy1Tdh
C3aQ5QmHHbCPYKeCOVQ4FZXEaOq3KV1lNeiH2KuKphuFbVIWquglYYfEBwRvuC0t
su2LnOyJWxb2nHZs9/2lHSWZJZAebU7b6LSZJtD3eS6jQV+X4MzROCG6FtUMLjS6
FaeQrCAF+wO3D67z6XAytLLNAo6Qqq9GiEVdrNJbSs1reo+4Y9NPqrjE0FbiFy7a
W+i6dZIaibqsycuqkTpLy95yIZYl82eh2wCC0uD3Pa/Sjjih+RRN99dR3hNNAsF9
Bfo0pO5B74O8e1Dynje9BD+RGI0LZ11tUjT8AS+e6f89vkNn6CeelOpNvbAjVH/Z
XHeza9DIfZ27FJYEXFuZ9sDYg1bP3/A6wmDxpOsm02HrAxKzQRt1iBwstgktlYLN
QqIMULYYVJjNhcDLJXayRCUVtorBoAlZCulQKHUkBrDzn7PdfkBlLt4xZg66uIyq
KTLQAacdmRXw54KC98g+jjPT0VgpayWBToUKXBVMC4hAxUWk+Dp+Klr2mW3+rbwD
JyVWEKhuZysFf1uSdYbZQSuoXsfXcjnM7AFQTbG7PTDOep7tOCPoGlLiQDE9wvSM
Eg7NmIwNV0J/G5WZUsnr5N2g+iUUM1NuTxO1LQbqCwZUagL75+vyDW+322FHkIjj
ZZuYHkeOzL3+4aSDBve6F/Au0PXISLa9E6k6abbsicyIbrHW7du1iSHubGpoWMTH
GiHiuni26Zv7oCTMXcig3r8Y/fF73F2p7V6d72M2TApqX0cbkuxEObqRCxyDVC8g
XTTqRfEpEjM6uMcZ0BFMnnayQWXZ7f5bFKsuqJyl/qg85kxZHgsV4bL6xfoIxdZX
AUGvbSx92WcUs29eSI82xbXQhwk1+Gxm4PeSMaJRNPmHjfnHhhNyYrAmQdxjmWG1
0ODesD2axxmcm+tLkUf32kyHoCqwHV+1MJ/XIHl0auoi6/jAhd5je5Khg9f1mjan
EEtI+HuNc5IIghCxM9rJHD0gDjGvuIlQx9TpkAYJiI2pAfx2nMbJL4BeJoGkoWvG
BK7drbnTvn+6UuXvH2H7ZifUdl1RapO8dhKEQb3Hnq2ZhZM4LPi4JyZEd4buMrTa
LpeeZ5BAyXLq6tCxvP7NwMYeyypyqptJStpW2PWSewz1B81CyDuhTbzfl3J7q7rZ
VPaq6usCpDq4KYyO4Fk66J+RTWNRDDpBg7c4v7Wb3dcIjknV/8XnWQZflm53ExWj
sxig8Cwnd7FZ8IcAiN4H7Wz3MOH7GF4LefCcnD1I9N79dUqZo7gBftht4iJH90U3
XaETuvZgl2hR3JNXoRulnHKqp6EozKO3STsOTiaiDeFzDSpJTp+ah0r2vEAslcEI
AC08Bm8J87i5P5nmFF/7DUiOEt0kqkaOmisntIdh8Gat+oqroilzDLTiFslw3xoZ
wMjihr5iba2iycdD65ytGHp5T2c0x8Va+Pi8Kom68rXtoHtFb/ZP8VWKtCsX3ZbK
3Llniv8kA4vrqqQfA0ZrSU2pGgl3uDOZ4nKZWQW6oAW7lM7/ePe0TXGiOJOyoPk+
Qr+2ZEMWJQsqvJG/bOOenaGHEJwXehoYtFfo+I1wRtf+gMwLDvKbZZrfefS1zhKE
o9DypHnQA4N4exdNiLJN4nj/40H6VUf+LUqruo9s1uNzuBcM3fe+SeGbC5LrteXC
FZWgWD6oZuh0appsxkAJV8IGjEvS8QxfGQ+v5P6bXsch2MyDutuV4NsmRiM6b7rd
OaRMEZL6hVjDrHoiLaZPAKJABxs8Dtmiy7uH9EWPMxE5z9Hm/qEnbqNvKZEXZp+7
pwTg9H6zbheOBXOz4QYIPuxj2u+Bst5wiN5A3kHu2VVsjfcGfknRMn8QeRdPvNVa
RFw0wK92ChxMhyEzuE54SGAB05/g2q5U0J4/19ST9P4bJORGUn1b+duVoJb5f/nJ
xBeCm/4ZDo+jFTFmyAWO2WZuC1HFtzD7+qqxO9SJxW3MFCZDw/H9O1473TgO4UFV
1oBEDbcKLJh8wjmyrEKKCKlm3cbzEYB4vL4XRvyavjS70zMzGTH8psvWLZVBHTYO
ZF2L/Hm4SzKIrbQ2/ZU/TS7leE/o8nhWo37DIINHfaSCG5CU8nx1yUZh/uQS7xLU
/irX69T6RgvUOjQoe6anqrFirRXIAaHYeJJOZyfFFsY4AqwyHVqlUHPUm124gWul
1sSHjifbD9K5Jw/vkZNLl7VmkZFoctFR0WtKW0/f+GVvw/a/5vABbK0ZjcRffLZs
S/0pMjGYzjxGQOzatthuuoadyzWNqC6H+R1TEsEME53vqblGZ75x8KNZqIdr9E/i
Q6Po7TMFknDMxXoNatabBgBxHQKQdjPJPphg3mRUVWeTaQFf/oQi1QeG1wLBruhw
GZPH9lgRWNE8wSCfmVlFK2FkpNolgYpJIHJWitk9DBK9gloTMApmL/PWldoZ8j++
XX7jrEi6woO2l8sFNQE62xOHJ6Len+7MJoK6O8RVKFuTolIDOc8sLYtvwGXGfSSo
j5AmikHJcpox0PWdnejdHyFBKX/Cgqg9uAuKLLLOSTR1GgdQIYZkT6JCTFs565oj
5F+0Qzqrx49vjekVPH/guPSDIUZY1+yKg9/mLtGP2M+4nM4c1MTRUbbRVswdR93h
xHS1IkRvVOZCSpSawoNUu53JK4g0JRsUuzK4GXoA7kldFUCNYeV7+6xHDQ3eiSJW
2z12YKwCbz3vqKGOS0Gcw1NlBe57Y6lBfMHcsn7gmnEu4UVZR19xgQHqGW78fxh6
GikLWkN2pPwzBu2hxY9Q7Hz5fAX5aPrvpP52WtMjNCFEreM3/5o4ubN0CwOzl5WV
WUoCU8RPBaBXXGJQWfiNyI3CbbGZ0RxCfH5n5U6BjI6H+hDuJzTmm/3lFauP7ojy
8BcuKEBHU2aeS4oSWSgR6nzWYoWnaj/oYDI1p03dZDh+ZLDAeZ9WZ3JuXlHw680b
rhGxPjB2TBs976AtMj66Vzq0nrvjPTkg4Lcz2X8oBscs1gmXbaaD6k/PmpWgPngL
Sxk+JVcAVNnNNQle2up2PyZg2o1AV+rf9A4SaSPlKl5/VisDyilM9dpVFxDUBxnt
3CCLjvDhjeFhrkgDSzfEbgv0S5n1gPoDYBhiOZMfOTg/PoW0hjxMypDB6AHamgdU
tTZdq0JFVdAKg72trjwEmv1Nz4mHlDnaD7NNs2kSvjAZeE3yn8gjUbMzuvmFNjpY
LHGORELkgZfy8QuMXDOJ9jzPWXUTaVffwi8i0vViDREOnl3Auqagwv8C8xCIwJW/
AXn7vVG3xQo5caWWZkFetS6gDaFl5T6T+ivD/dK7wcwUGkqlhbDj0WTdeHgtCaDN
Gkcf0mS+7pD/ioGKpoX3qVsMYoy45qGeityfFb/NcuSJHcm3DAyhqTze9FezHXAw
KBlOgMPntLki5HYSsG0dYK58ZUfPGDduFTI8yZ5r4eg7g54NFq9zukwwKgjzCYIt
DrnI2/OktqU9CTq6OHcutKVLX2ZxSJL9OHO+GKjPIqGm0kEXT7iM9N7f6F3Gfx5K
9OONzmEXjryTSvoNQ2C1oweAGHSSvOcpqKoy751lUH6comtPakp6GAW0wE61KHjx
SHBL8VKYpYc4SdD2/w+w/GCWzYShYUEpuvgCXOxi6AxRxlYFw+qxu6mnLucm/Qxz
4DNupysxS59vkeKNBMbxXIKXginyJvBMd/cM298MH9fz+gH6iQ+eyUUNzT+L7Mb/
+C0+PtqjOdJuHzZ1bfN7Z2bQwYIR1rdNhzi+NimRV/o25NAvxG0WiOHi8QRI5bDM
30IwenEwgyP7FYo06As7ntTogH8MzX2MFcjyB4qce0uL8RAt4cfqgAxez68Z4o4z
nsKmY3iUbUNXWeQsuySmfjX3hhiVjZhbng0InkCzZWpwdry8Pk394BJx7LrZnEU9
HrWBCFky1HgXuNTO7huMz5ixceGlZ0zqAVXbF7OdaCBpWOD75RubheumoDg+F7s2
DCGAVBtxJ6KHUGdMnRNbI+hL0HSEn69FLQqdPIEHNI9AgJ83j/Ad+Y+7NeIDqjei
9R4JjKoBLr+QMkKOwe+DCbf9Hnjo6NeMrvGvBrlrimoY7WT/HgzM0JiPplFtdgOl
zMdAQXAOm04jQDXlg6EBgizia8qbWL7/mU5iYrn9MlHZEacCqaYsDjNx5evTwGQj
IXEIho1au0Kud6vdT77NtXzWEQ6kHfwAqbgk8CIPS+cZZYHXyb4mNBAZ/Bys9lRk
uwXVBe2ZGXRdO23fyiDc2SVUHQH1tY/GMTMTpzZCXwAJ8mD5GcXlOcEM9K/8NA8a
m6vrI4tfQHD6sQCb3SVXVymyULrBGFj4D04vytpVRcF2P3ZWcTBxkXDB+WRuN9Gn
RjEwuEQLB4oCKXukoKIWezJfoGx0WLCABHW3wjvnVIx9spvSDARE09hrSEc8Wtog
jCMTQmKIjfQ7K5pCvd+zPmNkz0pNC0h7k+tItOhSrb6+NI583H4GExXYJ7aZKYOD
fZuAEVajt7nI16GXw7peplnN+XT4HSSqu+Q2KGfEgfIJYn1SUjqBIGHWQ1Pa3eR1
7lH77T1PS4Rb+HXRY8tPwEepfjsdoSyHFUqeNkwYniIrCrD0erYNr/QZfBfZhqzA
hfxkppvu9MyfUsRjl7PzhBmhV73koaWr716T2PMp/LxFx248jPdYSpY6qhg+3xHh
0+SHCEhGrh8yj3GNkjFyZEJscCYe1kbNBiErqF98AuhzNUkiODyIsqdXIuZZYOSt
gxQDhjdX6DPeHJQ04ZkNvte8Pwxw2VpINbfTXUoEwKXiR5rk/y+wZEPj/ArOdmXG
kZGczXVL7J/MYEH/xL3Bd64W8a4fKuHazQhVsfTjbAODtI5+a9yWUEyFWfEc0LyY
zQ1sNs60bqWhs4TnPFZhaasr76RZNht2nYdONb1I8WtbvaXjCqU2d8ce+1EDtwSL
clRWKXi85pT2Ki/9glVQNbiOz+1toOlyR/vNqATkrN5qXTzcItJ0OaqZ/sp9gtCn
PXPSmFr1YEHlYgSuhorexhsNE9I3cnWRnluTADCXzLog4kvqeCtIOoc43Edu8RGM
g1rWCsfpVUvx6BatV9ps+sOAcL+FiAFvSYLGSnIH+BepQqCSOXSZjhb1lMy5ed80
m2lpkjGjxYK149TEUOUbV1rZbkxKMUH826SoS5kx9RN8MoRI7BuLUqRGymEoRVGw
9iDceMyqJydV1dff0kaNYwdVDntL0yt5mfUyzEMKMmucoGjBXT4HGvOPkSKXyaTQ
ktMZxGx9EagwnjwFKu2GjFnUyos9oo4NLaCFYHxJQiN0uyu0OlEbz2TL3Ss1Fxc3
6Qtks/eZyC6A/UVRX8LvT6S4lXCJR5nVmD0bcBhs69yCkL0JsLJSEBsBAuFKKha4
uqI9iGmMBhdB27kMJta47t7oQ+iYF+nR9IzmzD9cTGizT5PZGZYr2fJHGWNVCkEZ
8e996V1MctMEdlMWFYvoZFSrUIv3jTTEY94AlbwbS6S4KnkQiISdAxJzvwxZytqO
zfRLaoKrt77t1r/8DLRmxT0VuHldEalpJxSPs5axVu/Lm8n4w8dPBAoCv4cwVl/c
o94ugeQnc/OvOiBOz+qu41aeSH7hClRfBvkGC2UyNeT8GnYusLATpSsEA62btpDu
41IcYHkQV1IhQkUezd/44AgZFloKUeba2dgsol0/zKD6nEEPEu/DfBRQ0q3rwWq4
n1km0Y8dTNO03mjKHz2Lu3guNdet+nGTZgKaFWBadma9dM0F15kgHpAPMXG1HVSs
A3X1xxgzP2x//bwF0h+vwdwpMlNRG04xsH7vi/hBMXSU/QYgcm27mjcHxaB3w+XY
Tnb1ut7cXc3lLdJ0k5wbsF9wpcDL/P/KzThtC4ARFMI0V9JM3MNXFZAgPdHVwcL8
jWq3rNhTfVZYEDrNUyrIHsj+7hYPf1DrjmyuqA2eykfQNjx4QiJk8BbyQGeyc13v
OsZxn8+XvHBRcodquylGi3idTcsg3Q2LHNG6DA4ew030tRpC1eOjUOdWkfA4ziUE
CeB+gVgEgc0Fwedm5+zy3a5evFHaHLeiDI6xdrvujSfTtyKVFN58sF2wnyLzXnY3
0D83G39BvxI4PQT0qpJMydOEfwqqaSb71KA+QqOx26s/xmYFVge0NNIAL28AXntY
YdF/eVJSsU7GKdd2SeeT+M+Kb9WttnJ4da7T0/PqSjYR24LZkkewV+LRwgIPfZrv
ofKql3qwgg672BBrjPZH6wT8dj50M1Qh6hRT8sRKhA1K3UxI9CYb/uw7QO+FxXLH
V7oVZKDgS/AJLqvqXXe9DCFxgf3BNIdMDkQg8Q+sFVyFzJd87B1wk8h+2XAQOc0f
M3n7ehz0ePQQemfvmlOCnZWFCMimJHIzKaSUxd+CLubxEtqJhRuhFF86ALT9tMrC
QCEUSrveQxmqVlPoCEdsFymHVw8GBx1CVQZyXKLzBzSWij4YfyNR7VjKthSu40oN
0spLVttUKpotus4/VMd9DNkMlN4JdnzCVkqriEOvIDuqXsHPnR/cuijIBvd4UZ6i
PFemKS0C/CmzUP2AXQcH73FJGmPUO/9T0OKTEItud8NGK+KTiVBcMKIgBc3b7XAV
JpfJPS5S7Zeg2Wz2kf0ADC+SL2IWbC0UiC0SIDaES1g/6pRnMSVd+oplZ8yZ6x2W
sOEnVQ2HTUKfKWPE3A3kmHUnT+AJ+0TBfU3EC3DHypr9qRim0Y9Kja3Vlh8w1erH
evxrhWvbg7K6GA8fJxkdcIHIrFCGUwT5+Ce4JpwO09fdgIRKlALQKPDgjvlDh0A7
XnDng2iDmgGCKvs1TOP2EhdxVOf8KjqsiG1RNqfhp81AKRjmBO4fau42wVPSVouc
GquckjNJ/OUWL4TRvK7Vys6/6zNcFlsFbtDaXGmvtHIQJmefdDFSm2d49gyZnNkV
axYB/QcYPZpZ5WgMJOY4nnLZWWQI8qC4cBOs8G2SjfDA2lb/h4x/EWy7PjAMLQbb
y1ZyItBiHrx40r9Tamb7lGbFi0npheB5WX/d3gp8nbhgGFQx3qDjlFrY7N1yna9o
DbIX25Fb0fzh7t7g6WpX6ysnGDEVilsxO44mj2Dk2Mt1mxLfdZOD4wYl8yYQnkFT
MPrKK/lctEH6Cq6kkuYhPq6mSCidZqlVlxhNDOhBuymhc6NqTb2FWgRFMK2tcqIw
TNLfOwrf4vx7VZ/ElAw3ggnUakzk+r5Y5a0vMnUcgu+khohLQ1xRe6tEKIcA7m9q
TKnGBboLyjMPwr1sBGcIXgzlykW1R5fUzWINdk7Jp9OsBloCFJBfk//+DgGOlhBx
ycW57FmAYaYTxLvTXhEpCpHX9J5RIF8TIIJr1RIIoU5JxG5Z0ivNwmHOFC0z1BL1
44bfZlDbjYgUTHq9Y1V4fsRoThcoktVMI/csYNuNKdcb3o2Jpm4C7H09agd6qYtw
5PKnulMkPQM1rQl6AceGO1N6nD36B1Zj7+4Un1vgUz6drBQrtZ8zIeHliDPzyxLE
Vz0ze+QH0f3GyY23R/V44WSz/OdmlJ0lGEX6wGB6ZCam5CIP6YzD+NOTGTqMW1wr
GBTWwfnynT2MdadozxZFjjc5h/2hFWms26Z3OZGfw7MjMsCZyBj/Z8SdF5qPVgSy
HALsTrWwulg+N8Nin4+IoYdf3nnGbQX8ANnbYD/Yg7UaE6rZVg0FuqutFU1ju8ZG
cxx1T1tr5aoQlPkhUNEsR+V7P83d0gvSRQiuatc5EhmXIA3C+CGiYseltOz3uOvi
SGVBwW8YRaDD63+McqzKPbgpkczAfHZhRqVDyXCA3aWe4t/egKVnQeIRADTPt8hS
XZsTJDA2AEfVOwOe3mQ6OyrT+iPp41pZQWoGruQwKx8+HuGYfra9zZWrlatDvdq6
MX5t7mo1VOo+/xTRFf/V3QtYlSJthBjNunZAPFyP7P40jLJP7ZcAcYgkZiIagL2Q
7IUlpIosqo4tROYtAHlaV9YrmtWhBnb/6pKImxURGf+OpfUHCY3esLaoOwgWWxSE
b3XedSuVR2OLWOn28F/OYCHq37e+bua+zsu4LLcULVBFjeDOEWmBI/MzsAfVxvkV
1UhYqedpfGnzhkIJiaCqqQAuhTdNKTi5fvHlqwQbfZWJDEQlv+SIoDMqq9x7yvqp
akdOsZCzJ2zbx8FdWEZwpJxx+cr4CQOpYPHNvkXz6ZpyGuI+yO7evaxOiTZt/dcu
L0QuhEpCHNMPwukMLIA4KXNRDMHlJiESu+jS5sAFwuT+UXSeZo5MszwIwqvYZoKD
G6NiEAvd6zlwhj7KuVI6lx5+TRfoRu85SE3WUM0ZF4GQrew58BAczomGkfnUTwqP
8wM/QIQl4+xGiEI5cdgs/Lwh36q1DKOPTbvmporkQm2t/i3UWrsTX6C9PZS08wMW
Xx3Blv64m+uZ4usWo9vEF2Jwx8AK0EavXc22AmhUE5dePSnNCZUxvcLPPsAyjoaB
A8rHwc+wJngKcsCGueh7B1/ONEh8uh0LwXiJ3sil4WKrAelM7z5F9AsJU8RiYFKB
5b7oDU6eogFQvCHig43Bbjl5VksuAHeZttEKA2dKsC6s6uVcD14DNdgQ345CgFle
8+GwcY/G+9u46rfISUwDrfYuAhpmlKh8OB6qPQ2jNfr7dkVNac1Ta3cDQTbyp31X
fHCJA2trEl7CVSKBH+nhSds1CoU2VuCgiRQY0c9nxzWGjzBLeLzw9S1/X0nOQlkC
1T8BZ9PD1GbCQoy0u+kuLUI3xMnr8xs3ZlU0twiZZCTtfF2+tmH0GlWeBFMnuiuS
mKzYC9Svewj3vHKNop5chYUFYc2GgawKCvKGXJcvHxincIEAa59GXohG0SYHOy/X
/6QnSKqnd+keOmMGr3QFNd2rUykm7mwD/80YaWvY1v42XAJ1NtL0IPsunbG3HcjV
o+wICaChU4kBM9U0gPtcDINetTnMMg6ZBG+sGd20/NyWVXMa2vGGaD91N/yYSuRF
EB2umrcBORsFsUDmK3RDej2hSSKkbkHIePuavXH77c6uaBGM+ZCz4MaNZZ5FMXrs
TgZhzlXZ02/ZLAdk05cQcwEBd5rvB8U0/XJTsMeOSevNyaXXMZE6bkQjPfyeIQiJ
AoRJ5dRXFvj0Va1JnOBmNiA4u93m1bXQwEBfLkmtyQvlQbGcVYVySh8CKhIoYI0J
/WEdwptPhS7Nz2OH4NNRihevSdtXCg+K1+aZ3InmT1XhNkHjL3q8niAfJaojrgSS
Vj+1pEMBqj663pKSc2wvX8EHhKVg0yGwl20NS5UngTygpI88DJi8kfu2fppuSCFz
LwjbMuaIHAi7pZdEOnkcoONilmxAL52FMXMOYOdJWHbt4i3FcckTBibjReZ3b7yG
zKrfR/yRH/Ov6kuPGbGQCiH6/h1rb5ud9ELJSBNUwDhLbJqD0m4/MUkU4wurNVCQ
o5EPonesO6+m4nAEJZFKDUqE87IIPi4M5sYHTfqLFZcDCLZnuobso5TljGa9ibfX
8oisDgX/JIF4WC8kncPybGlfi4sqa8KAkTAX1Kt3MdPIXZVKttuhcceEznS2rkKf
H3mYyTX3Xt7DoanNqDoWGXfvXpYyALb0z1cyEOwNamb+/mrnsniPnojGACosnH3a
OlQYQWTG8nbD76pWQg1oicaLY42tVL2RLaMJOnVbvhjxkWd4PJTTWzxaJBJOnAx5
VUDxwMJrAvtm77BFtUzHtF4CtyXM4n4fMIwsFdvKpg2PsIKz98lG1+2uhaj//ZRc
R4pjz3Usjxk/+qvq6mULD8bIuJCsErnPjkXOWGuXV2FNqGRjNWJVLWpgMTYo+VJI
1spScBY3Bl2dIkTszyalm1MoXOiB3CYqvVwODXy82U+9b4MPA/hg/eQyUacsivGK
KqkyKi3uJz+PaSabKsHkpJ5+duVoG1GaqVMZSV99RGFEbJbDa4EHu+pTLW702RfV
/JSX0JSyUn3GOS7iL+aqjwd5R+r06O8Wno8VyX3/mYRCeg9/fDgERoo87AwsUpE8
ARpClqV0ZPmuyZgzx0Xw98MZaI3Ou6/IZheegxTFCthyh45RtRPVsOW2rAPjtTPq
MQjg9W6GtbaEQDv4nZ1efCvVpRyfXHMcIk/UmFOb9PUy/ERVdfohtUTaYPvaC8Gd
gW0jf8jcEyH+3XSYeiXCcd1fj9ph4xfpTbZI6UkNIRE1Q7MZQksEjyYp6mGxW4L6
s1gqFb4nzjd930EkgP4wbtHLlBr+SgWbDJ4DtLJ3UhzGK9/XrUXDtLXMuhqpGD3n
JewK8A0yqvHCYTnzj7LjiOGOn/TE7h2Vvp2WB5ivhpnQwRPofqKRWBDsxWDZAoKm
OjlwBZIY45ALGfP68SGncjeVGF1Bugc7KRaqfMnFY3MxdWWh2j2jYYg21vzVb8z5
WcI4Lc4S0YySsThblLbuNhX7zA9HiNqoOZCvSs6cH5/QLNr0rqExiEh88+GzW4uS
QFgE2tSVZfv7clKxLo39NDvhamknxKxs9GnuwPJRKNLYp2ieQE922mOAscPNf6iA
oaqBdF1Gu45N764H5WOBACBVjXd+zjYV4KhpH35B/1rctcZKFesIr4A1ioqT64Xy
aj6enHOV/kEc/M40hMfjhhGmW6G0dGKPOWXlBixSS4LRtoTJW5Y0INndxFFjCwvd
KlbupkyIfpEEh3Mneiejtc2cse1jr6esizIsB8GlrWIwVYQV1AfQDn/oCychulvc
frHvxw3bY7R4KjjqwPVvjfbgUNr2MlcI40QXpWag30fORGqgDLVcTV/4gp0SBVW/
uRs18agQfLHOYLWGIhJ9/n5NblQf8h7P9z5FWyg5AhKWa8z/Lrjg5+UdCaOIhaz3
9XNX6jiyzAHTQB+VVxUViK7XbzXhAJgA+FynX1FDZJi/+N1Ox3re1Pb662umc/Ig
NVqfCcCdM0LTaWS87dUMK3pYUTw1UteklgZX4Cnb73QYAHci9ad/e/tEP1yqWgKf
KDUcjcMylzNmeUd/vP04gJqgbasJgszOEbAg3+5WifCoj8vaZaXWAAJZkVpJsofn
iaxS/bdQecY+lZjBb6WkDGhdp4IYH4ZXn/IluhXeyfs4WYBpYwac7pjl9cQyVdXi
4FsSFTu7QAOSpUI0iTcLy/bnjMCsOTg4KgfWtB/wdRg3HB3bdh5ElGXYxWQ6os+b
B7083R59JHL38YsZZ4xONTMo4QhJIq2VrDZhhPgdcx6WFmi24z87glr7B17iAcvg
+EA0jQ/O4cx3L18X0Gjn0Nynpf2fDjLY4142YDssjgxXhlhwdxaKl7GXo0OdYdmI
tDMEe6/ylw0PKRBaTB1R9LE8IRioS6ICR3CX6MVrhhU8OIeKoktOVSaD8gHY7XO2
57UyfQ1+qfs2KjVdut2AV7spjwikk6wqT9Vv08N6sXkYiG9cTNzbxe6JK5bERuza
R7ALs785OE6NclgRMSpLOmU2xmJVM6qGQXZp7qI+CxpNy9W7Gksv18NLmJbB+IAi
3oRV78XFCQxhA8CIBeA/kKz+5jh13f9P85foCnAjtcMpzsBvp3zHgPCk5DJCYUSe
CUbfJIqId19iNOw6sRy1vLnjqq54xz75dhe6a4CfutFVY/Kv4CB7ZwgE9siK4oOu
et2T9UQRoF1g4EQpf/7OoLoqvcPtxp2a0mKRHA6sM3QSlucMx1UgQqRf7jOorge4
/jKAOkVDr7v11N3xahZ8QKjxPnw2WBONqF74KT0ZGEQ253wgt/KrQEE4kiMUDK5L
d6Y0UF6N8hI5CnyLka+Hm84nP43bSdATFz1sge5diKa3P3+qUtTbn61S1V8sfqRm
9dmW1c+vLJwRqnUif9wayVAa7v8KkkbZ2guwvpTXLR23hqSTYKEpjDzVIQ6iFNdz
tSWzqZm43GwGEmBHPLFYnyLeLBbM8NOr6HcEpmlg4koLyyWQf72LH7SK3Fg49VJe
/fkvjl4IjpcP8f9Gzftzz0othjpaxVq7Pk7gt9cNF/ES0q7jOw6RL0Z/SMoM6zCw
Fou5afZm+2kUJRonUW8/gvgbec+DiEJY7ZwJKnKiPCQ8PkBxnqzFs0Mbb1e1pR+H
iXBEMkdQoH9r0o4zBaYqce7C3wjvtZqslaBgu9fypW/7Xj6gU4MYryCurqm822O/
4vuKxoQB1nMx2qbQPNsXzx4lGILJ1M5uUrrQbfsheFFbzinMvr2/0JsCKlygN3Zk
qhLAejPySWxYwS3Enz/AQa9/AKlwxm15oK3wOmdX1U2f+lS0EnnR/VUoftfG9JnN
xD0zAW121ZiRunpZghl26Xq7qqDwWmhgeRx3L7tBCaiPQ9lcQg0xDUPX3s0ch+Wl
ASLxS8H85lPdbkLsKU3fgkEGLcWGtbWZM+DxVtzgkvyfNGn+V4hwWjTzM9tVAdHX
GYrbCP27NemKbAgmaNnvZnYZy3JhQ4RkEZp82qKU6Sr+cmdLCwq9CKkSMuVZsSbx
Xi69AdhuWet1LzA+R9AMwMEippeB6Gc7obGU0Kl7rdHufoJcgywBjOPPSatSgYbD
tbF7mftwgcLYpuiRlhrP8R8jmJBmMJjCiGIT+QvwtQTWaaaC270Gp2moNtGfm4Bp
e0QXjhwSCtW+ZrRzplZ0rbLq6eUTDJac2mpchtZcWQK+553XJSXiXs0zTq2Gj0FE
RCWA3ojHxWHNq/MqX96dLyGP6FGhgBeLOYT3XfMEaM0YkL8OlngeTb/3BCXnpaCW
m8KB8rtARuZBci1/0/Ia/tSI4fliJcXifwxjn5kp7fXJ+ByvHQXjP6w0+f8P63T4
2WY107tygAGCEuH1iYI3xTdqD9cMKIrHG//WpsCcaZPVtCgxZtueFlM8/r5xt05Z
FfdFSMQyMfFnY2FYjrn3iM1so2egOUd/AcmpeD+XCGn2CBn3GZtUvHgmVe9BjX1V
+4K67aksUOIc+Y2qPKa6EXWpSYtcHWiP1Bg4xbKuU5V9LkxfFes79dPGoaxNWkcD
Bz5yrNFOecpgUqRRPEtQBvymW7jd9u4FWA+NLY0QeMNZ2sLb0x0Lv31ZkMKTAW9y
2TmznE00Mp5hjeLLzbmopBD75LnzyOSrx2tlwofJEiISfjGr76rDDvVDWps9LSD3
UJ4MNiL3M+42rVgw6s3V7eMcj7iKkCltadH5USioFU/WAQ/+YiZ7xkX0D+IwkVrq
qQyVUBYwFno+kheRdBWsmcoZWFbdW0Xl+Quv3u3RaTt3YkA8XHnral2aOiNPcHtP
hVGRLj/TB+fh6o3UY4qfThKzYj8w/iICxRzUGgKPdrBywtQTbCJrrgpRoKmbzjTr
FSzOf7blKNzdP4TDXLj9WJAPFRd4CxXlhk5T/4mAbQaKul5xmlTkDp9vhlAHs2RZ
4VSgclqHAFeAsuw3t4DKN395u1aAAJAl2GNsE/oyxJiNcmAtGXD4fgShsV/aOqqC
0e4WMz05///zUmQQt4+Hbu9NVmRM6ei5mnxXzYaxa1G/zBSX1wr2JprrmuPsKWwh
9yZx0H2/+SkLrSWjYzCNi2XnGtjuBZ3uc8wMa3+e6kAYHDRkiJczU/psj2uY9C2K
LcwXn4/AbYCpUnMziW/90KCSwN+rQUmkgnah4SkWMUQIb3VBoKYiKKkwnv2RwZa7
n7gtUGNyEsAoEuzckXkEy0T9etWf5ng72Pyk1g6BzDOzVZwWX5USsF4tfmNMa4Es
s1FpeWK5n2aIXQ1OikHBuAOz8X3a/qbOHvMJZxL3uX58IyEH8+4mrYieH91QgZrH
BOM6qTJFh8yh2sTUpzEWs+PgbP7lz9tGAb789UlEMRIoeID9nQ4uBFvYv4wR+mnv
4WbDIDj91KBz21J5gPQxsOtu6qCHXtYX9QZ9t7KBx4VNaC5+hdk90Ma7C6yk9kJm
Ht4nZvowDrwZAQa2JTAR8Q9JW4RSMkCZ8BdpStWHM+X1QHNvlRbhSeMLC0WnqUrB
V1XhU/i3Y5cboi+UDtg+YubnwxdMV+R3JrVPNJlGeCeKNzzTLYM6hff/i2IGCJg6
V48XxEVSHUT2rFLOwvxYguTews/xh61bOyhpP7wDF9FcSAseU3Cb4nKycDo4I73c
5HypsKy9KftvbSEizhhuCrMDuHRPxB7dK774x8vASDMtA7k6UelikZyCHnv84rVm
sfZXit4WBO2d6EH6iOTwT20fzisUyjBmll0t4yAeF7wIArhbboPxBPE+CBa7qD6V
f4O2wq6YIW2ghvVx+vYX4X7fjAVammOswNvrUTsVMt4yxGNXF+h0nGm6e5sDiPks
lTlza+Atm6yyuwucIIPgvyWFWL62AKi0kVxRwJHbUZnd2SN0QffiLRieF1Gh3cT/
HdSCirjhsKeuarJWlUbjfg5xYhwML4QYJgasqvtzwpQIVw+591fJqWVRrp9IccrO
LArSY/BAJZnE+Qj75G1gukxxaQv3E9U4L55TsTZ60lGeQKUgLVt6Nh35pUfr+l13
dbuVyPj4w990lXzEj6cQC8BN7Wx5Nvp0XYM+Ko3yDEAeaNp8GhfkPO+44ODt/Adp
rQbrDTKVe5CfnL2gWNYeCclcgArmJOEElGxCjV+4goCVCziRIETcNifJ62HsVh7v
/VevCbzDs0sfHGqcSHWXAqkf/ocMDXUAgoSTNLE8hvHdzH//FFmO09s5YX0cl3vP
v7PxYP5o8NLvWDT2hINJL0De0g0UDHbQx6YckHgGBT96pyA+H/butERshyvM5p8Z
4wni/muOenlAKZA0gF+h4uSmR/lYso/IcKLlm0Khrhn2YO4TX4UE+wEV/wrOLf9i
UgjgyPqKeoGVr/86xyC7EFyYh4b6X77+5IavSeqFyDJXXX0yhk2mr9+/XzKmoovW
x3waCmAcUnzvaZ9Nl8dFnlLguP1Wj7FG5aZyEuPZGvO9Bhj2A7ObkZQaKPIWbWDy
zUn7QtsDZWT+6kRIIYt+5fbbZXOSOrsuvQpxF3cmR+IwEMg6xY2AkIAjzdgKGs0e
KmoLNLlgxT91ko5W8BAnEHnTdtU3PnRDFxZjCGQZualr60Q+aeuYqWbtXY5WmvBQ
gogL+Z/T+cWsFQrgOBSadU8fwKxt1vpY+PV6pLQMW5tAkzYbkIMM/y34jsmHKnyC
hTZ2evRRiwXjx3SO/3EqUeQde+W111sy8peY7iJo6FeQO8X5RsdeDwnNfQBLaTu4
0z72O8cXuZnL/3Z6WSoeFLS8tE+eIDtVZo5OBTxMb8CEb3FyZICIDdocRhwJtuE9
ESQqfCotPg/+ZsCRlfcx7UJ39ib8Eoe/pedEMLSwAUOhbEriVkMu3238uIA7iWBy
5FML/DwAxutD2bIjOcQVdWzArF5+v4WzcWfoMLiNjSaNyhyDilHm/gWaglerBBCU
LV5yfylUfHkz4GTZ7w2ZCk60O8b5h+v7V1l2k+pzLCc4FnZBpLOE0mLdVnjcvyIe
tME8z+qFE5arEBiROknwGc3KYKJom4ik8aglCzgko7ESdip/nLNVj6Cus9Q7ELVS
HE1l91MjsFLl/nStXlin245yiuTmWRoCKE8XEWPDyEU6a0uSjlJiOXxiEHCKVepQ
f/OX8729v8+j2326NKytI+J80svxFEzYj1f+VlY6QhkP73FgN9xgRTzMVNuXtgDB
psAnfVQjg2GPrYACaEwvqNVIhXuGmZmukgZLaTpQj5NpH7K6sYNJXv+H+VK794ri
1eJ/0AwJLySYiiHSHBu2U2xNbzThX6AAGakg7MMpLr8WIpqewAKuLnVIx47S/ZGw
TnaZkmAjuB7w0lyLm9YqhZDJV9iAKokb7G2D0SYUyPvwoOq4T4tNu0ORxAp2UKoR
SnNHGS36ykzKKjekrNCuP0SP3AQXshLLljEPXrarFRhBYSz0psrA6ac3Q6qNGEIu
TNd5NqNx2Zh9JJeYTqcThQ8Qq7MEZJDHAI0mvv7IVp1AcJAz9J7z1hYpPynhbmjB
L9tuOupyFjEe/dk6Y12HXjEQyWsoLJpB9T5O5vNhDpZTIfyWCcikfCUJq3kV9eYK
Bm/PaE5yDv9n4s8RxQohTmAAzTeEm948DBw+ZoU++HEpYU0+5ODcJ/mIIvwWaH1h
oJDEVwnyCRKVU1qz8xNaP0HKUilWXKvG9SrJt6vX+Ec1SHF5aMlanCzR7bxpWKR2
E6vYtvBptvIonkF93mB1uQZGda6hleC8q/zwZVpFY/sXOgfsORlRBdcA1JIUW6u1
y3koVDdvS1oUGjgrrW4KeQH1DytVyzFRg1lt+mAAUoDJELgMb1/BuYxsSy79dwWk
VwY0agusnuGTRoP207YDuhAjSmrdwiOuGp6zgNHEf06jM/E15ugonXLIKFkJ5/xQ
J3KjtP3epOiBv5tyORKpffd1jZRlBGUvceDM34dNIXjEdjSqxcK8fbspE/ArvsTP
ayjXctEBZBFtyvrUtFQo3tgG1esTMz1bh8KDixajCq8v8uxQSGzycUGX+IYFKCWy
X2JfiTktjOC0RNg09YlqvnRKlu7HCX78kmwe0qn6nQKDXlQF+2yWD3n7HLtmIDIH
HF1ev7lpLOofYg45mUjOZ3fcU+USfckerwUIbHcLnKzStot+2rzyeOwRv6TLvEwz
tI9tacJjFzklzQEt1PkIkpk7u0t6tDtQEuW7BRqI/H8VM5Xza9dMojMwoQ8bFaLD
v1SQHbYXS/v2ryYRbBBzmhlmHZ3oW9auyI1TsQjBoXUYUXt0FukOAZZLicBvtM1+
gNgxBIEbDXbdf/TdokLdV0nhf7QfAVIOoGvNhEvLGbRKhGya57rMTL4a2R3Ap8PQ
sPTYf03DMeqOoV4jLm7a753ynV9+S8Ddw/bK9wJy4U7Cm0EyFdmElcZDacBbrU3P
a6/oTmij19sWCl+Bv4y5CYyBQ/Q3/ublGGB4a+pDFYhkW18DkF1vVQkzvb+HVRY4
tkl/N3dy2qR22//kyNk/B00SBX4Dp/3A0Y3EBiyrQzmoiKNYbdww+v/E8FWkZoUD
/0QuqR+OkF1ZPa7Vsn1VOiYzc7T4M1DIMj5mj3g+8h180nt4ZICKE4ersdAEfqQ/
dtN0nv4OBKyB8NTOAYNLrj21WWQOqNVVtyUTZgO0gDrMOS8sghHKRiAUygA3RtFn
n6IT6nqm6yA7/LFYq+qPAk4oLKn/9fqRbEulGEav0nOaXkoFIzbZzPv1Hfx1isM5
M+1PIdZqCtzc9roKiPfnaaoYakTd6nH9FnZyQJ/BST1oILcbYh5t9RX30cOxXEhS
H34l4y3J2y7gZxLN/+k+j0xc13j5XAfMznH94luUvlVaHcLIL39fuU6/t9fAwOsp
kCQ4ndemn+TlB1cRHoBC0TuxfCAavDzqrn8qG70cy4dszMEHGqe2yO//4Rbf5JHa
`pragma protect end_protected
