`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OVSojrQzQiK+owY4MJcc1Fycx+/Ajc+QElIl3ZSSS9Vniyr+artolbHz8e7ego0Q
3fm9Rm4UyxrkZUulvV3tYluXdvlLx6lloBq4ZX0Vpuc8xp6FqEc44K5ONC1XjDkd
nAJ6p5zTrA11oxQUJjkyQi/2oqXVaGMw7oi0hFjEQGg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14112)
4+BlKXiJEgicruOcoZWiodH2o3FWUr3JdAnkMsb2EmPRwT6CVUGqQJzX+GzTRoHF
ibYhBQmUs55KChvvskg/LbK0OOxg5kzfhStl6sYysjTzrZ9FSGcqGPQNXEJBykex
+A/NC0d3A8W5nDPLVLiPbyF1WXjp2anubSk8vvkXyhBjrJYUXERm6v4yhEOqB6nU
0eikaERmyjMThjyFkTNUrIDeFLhWT10cJS+7JyeRFAAwLq+8PkldzrJ/DSeqyao/
3GiZjlrg1xMMR9nGZ35ndDe588kX+U+uPqh3aW0xPjogeqgbJeY4UKYj0EV8Yl0a
neMWmavFM2cGRcD6zeuNYWXREXPjugGVSWFv1oa44ZrDZrpIbVy7ABkViMh5Aqwo
n9J0/aCk41+VUud6cCtMChV58J6LwBDCaf0yt4CpCYk758gKu42e7fw2ZdfYVfi9
IubkPkUVTTlHyK3YLS3F03Vs+oq8SjHfWQlfOAcNstQTrC9LhD6629NEG99tHnii
9yEeDAUekuJJXQl3PaC1JV9eCzLO68/rjGjwf8LwiHZxlXKECXVnetvwjbzc6UTR
PIOZ6NJ6uEtNpx8RxmlSMRkAJGgKKPDmiXWfAmVRnvnqi3WpgVHQVmxj2XgLaJQ3
7NTxQ2vFOLRrJczZ9mPCOCsNR0TCND7iYosB3X/1gQPpYENI+apS7Id3j11q0/AW
L02M3vhxsLEtLEXSoQhFJIeChuILxGVpHcRT5s0/1i693prKhWvlstVVxHarTo8U
Et2y9XIjmo9YeggLzWOz/okZxGRBlN6KZj2IHlU3JvzMZmiwxLQFR5w2NPxHeSH0
WgFgM/dwICVRfgDqboVZVoPwnQKY64mvejBqORcv+C5YgR26DXGDThRFtLO3Tj/H
y6mQEA+Fk/KVDMeBHEBBf1u7qBMrc23GeOXXtyZqx/WOFq6XmlbdWp/cC/7efEk+
m1C+eAhQ3DaPkmMFA1X2e43osK2Natno4AGMaN/S2im979t9GrzGVaafHymXWt0f
YddO0gbJQqUyM7IoT4d4PLYyigpHFvrcUVu1Ltg4nCq90y05b39t6lusAc6sYiyY
8lfk5YyyGU417trY1HBqXOwsQ4qg9N9tpCSLBDiWpcEaWwi397u8L+LKMFk/MDGT
1LvTf7KXKg4YTdm8bOMYEDWgP/a2h56gB/0QiQSMI/thyyFDhp6qP5cJprbKwC65
4o9fp4lwybplKfQn5HpwWELzfsQ1iTPkapP/28WYY9kXye10YFQQVIlsTyUugZfe
dRhbR0q8zEnY/OViNS6Rr0k3TVOlpVod4i8Ol8WtHB8YJkc8luFR1JCNu4cpQEZz
OTY7y10q10w8uNSgEsKDjtlhdisGR1WRn8gtgX07EKJwMP1llJZOds3qdpY+eoBX
5+W9YuSk4FUyZBXCX+M0aOSlHSnnCfMzWtH/W8IkVb6VPTb/FCRIihKNhPWMBPK7
5mt9zNObHBs4LM0uvupBE7etTZQwjayFFXrQGohSi/j+AU5qKc6PqmKNN57Zki+B
oInfJJh8wuin4i7M2GDeh9iJD4zgWgtLoN9zG7jLggbr18hI9Nx0uT0o+3cVutK6
rPGg3bBSJBk5V/29NznJIqYAjzL5Fmb0xGiKwuMvvoVma7f35o9Vvd8trF1qXsze
fq8AlCMrMGLmW+RRrteMSQWHJvCRv3FMf8BYAV6croaWQJWSzz0QyqCxxuacScN9
cSSpHy+A0+nhTxcGvx7Q80MShAJElCFPoL/w53Aug7imQshTqd3YL7Sk0ijOg7ju
G7oL7TRUq6WhNoTuIuQsFSiK5T0P8c169PxJejPqnVD4VU4osJD9axR3mPUSBmPn
16UrN21V8WvM2yfMPUzLwI7Bm1Al8uVHgPBQrR1ZSFLLtL0gGgjSRnxbpx6fNaY6
s139mmlNthbEtUz5JgHkOEddTs1vbCNV/QjNuqOxH0erSW+oWPD4DIskLabENl7X
yj1ZkUpu5GgOaZrQmtIboBD1aVTqr6vUdbjRnLNN49l1oRU2bKXbO60Ky9X3M0Nf
4ejCpfZSJQw/r9Kav9yHsf/4/AMDXT7rXDzm8/2HsjYiSsaVRKkfpOlfYWTkn4N2
x6BpWSSIP1goxjR+8T2vMJmOXJ+8UeIjoC+lOwY9ZofKoQF3y6QwZHaYq3QEmH2N
uHfHTNMbm/6q9QxEI3qLRN7ww8plytaHrsTTF2tEkUHkmj97gOEi3MciE2/SJ8Sv
mqCdIHiIfq5I2HDo20yTaBVySruspHUv6M60KGCJGUncgJkPM4ZXdGVnwpBoYYI+
Sr2DA1UXi+SbyplfyXY7XkQ8R+mJFCTrTUCy7TCTqcOClYmR/2U2DvZyqKtBnDMr
0K85Bfq0TSRsyYotJZdbQOR8KQwyyd7y19nnTdkS6v+ojDl3HsJeC4qOD7YXSTMC
WDiHkXYVI/v5tBk+wfIwPlGviRQ3mHaYjUy/boUiWy4Pj4YAKPughQT15OjgnE6z
CBOuwxdk0RxqDhyRGapquwQB98JUvyLPL/Yz0j6KVxK4nWuPv/v5itU36YHmGDja
z0oLsjbLhdryxFCxnmOFl1fmRbtgw2VoNLgjmDru4tJ/M7iPph0sdb+KNqImGZXa
O3nX9cyV4/QK19G8CY/ocAZItYzDzrsTLgYFoD5HJVY2QpBzpCduKJTYsQ7hVNZH
Gs1E21kN9Ogs5z8dn6lql34wzCMEE1rVMb25jMlXyW2tBjCDljwLoox2SEjxNBA0
X6Mtv7BQjffKDQ+h/0cvAgPAWSb4VeJ/hj9q46k60eG5o49uZBso9pH2y2R9gyl5
R7I4xqKnQagcA49snCzmIZ5QIOqyEFl2uIFE36SWpepw9JPddx0IICHP5229bY8l
AbeDNwCMhEjmXxDhCGpptUl1l5d1oUX8tmnXscbV+i2jQZi0gqgoDpzmQaKCreSp
FpLIxT6+cTkvk4/k9/7QrW6RAOXT1fUt3v6ZAS07O/UsVLgIdwf0PzvtsXh0DftF
U+pnc7XrYXyb4OMs6oRPiprOmSOgkSLd0dB6QRjQu41FUeY1g11j+cWx3YtW64dB
xTwDVwWKvnDWW9jubi2Ks/8JRrK3XSpDU4l8hfZdHZVsMWND6KMuyE1G3872gEnP
LkACdvr4e6H/ZVqJTwVq7oZfuwj7PQtd365i29TIx6BenwgI1uiv+vPF+cID6AGg
igUsbxwq3opAOb8j1TlfIlSHT4CLHHEtrbWI7SVPK++xLVP3OU0uzUXqM0qEVLMJ
12h1skr3mO/VcKaWNbDqSQGqZhLWY4m5wre4Cc7smGgqbgGcagl96eis1LdUxv1R
TyjtbLUJtT2C5g8k+eIQ8CPYe0aX5PoKSw8G14jlNOeDkALt6FY2VcapZAzfTzGc
bzP3fTPkxmDdDaNK5tw9/EiYwWcV9i14AHKuvC7BJ4DB8UuptqvHFh2x5GCmQro3
RuE/kPkNZ2aVEgQ6C2aSA2K6xBe/z6ehgrdLVPDnerVrrbR0RDa+5dj3OGbNwr/g
OqoDlfKq5rSCsrVN7gt1cOfQ2E+YXhmkBM/3tOZubatLN9GdseIQY7YpsWkfGFXk
3UpRzj+MFh7++D7R/qXNPc0g+mkfsHyUy+iKz/P73426ZdXT6d1YlddjJD/lvaVV
iqctXqmm9ph7Lz+8VpgOiKfRCOg0oBKg/aR/lBd2TvI6oKwW2mh7ofpOAkxVaMEk
92Xt8/530a1jzh7PwCRGMA3qkWkjO/yGBOGKAWSH367j4pUR1JDUF1qnEyhDNZCV
+Hqv0//zfKFm6G6cdKQQbzxbObTJDvti+0jS+if5KQSm70/VnM7ItQC71JcfJdq1
evE6non9Gi3mwmq0qGbfcvVCMArK1UQYPcHX5RcSG45m5OIxUcLamLL4kVVCMDTD
ZB2Y2bZzpvmHLa5hQmWbt9kxDxZJRX9qb7NDLE5mrsywbeoQz+6QVAtxZqwNVvmq
SsxlTZhu1Z0PLn8ARxjYiJax6pBA0KDiw6xVAwMIHJOs+ApZpAHUCgP//hIdnQAc
tgGCQhSuF1tTrMjgisQhFC/xV900iTf/TVq0wTZJtg5sfCEN9EmKlAETh5b7fqb+
ur4OYYfd0RYANUuFdepKZt6FaNKFQ7hq7iRsicolKDa8kEf+bAUHtvXIp0xqGx+/
QUTFKDSgfj/dVYjCmp0RzxmqLb0NqL1kR4hbCFTYlJscJPJj8lJC9A9bb76vwRJk
Vz03du9tTNMtOEdYqUs8kT3W7QwgPWySbMSqjnYlersv4IvxMpl20HETWTWheCJo
hck2RNWa4GsYs2UMEK18pvsOq7kuLV49aV50DWshMiTpoJfpzJgmKmjnw+5BJrHx
nCFOcUm/G6bSQpY9NUmDWi6hos2AeSPJmNTaLHYnq81Y3Ko7WLHTDNGzkzP04umi
BMANJ77CmZaGQjAld1DjYBEHMe1PCc8DD0v3lpfvEEnL8NKyZeCwJ2xB/oIdr/28
QL9r5D3/1uJUK1oc6PnpZU/opMJqLoh1oevmzfx/v+BsmmWxnXgyQa3phYgF0LXe
o9yLeqRnzowibo51UuRhH1m973g4xvDOGeH9kbR2MS48WyXQpHIO9iW1KijSaXW+
7Hcrsgia4cu7Y9HCBiU6lo//4AfppzbAhQVAxzgJsgL0qAGqkvAMGgWdDaz4S5Ey
cPhoGJyoOCNlmo0EPpwVRK7KnjzkFt8Rk7yU6qv34BioRcSj0wphsJs0r8ubddya
ySfrSQhxY7uQ9HhWOfrDwPMhc7GhqViZUr7a8Pw7pM0dmZFqz0WOwPzaiQTi9X/A
Gp+Q53Suk248pDi3SZAW9u17cOxB3yqS3eVQrUUr0vH3vJSOVwMIC1qoX5ClVdyX
0CbR3h2O50i/NSdNjrQdy0b651klpRZxyLK3nGu1/YlSscHbTuplAAO37CTU4hQD
VhzbXYmY0Nxg2WdF83dar9CR+7fvmtVGEyM+GvrKAjGFh9P9+WtMzcSzQxumHhII
NQOAg7V3S6Z+xfEQcvDYM5CJX/PkdL1L0a0ToGDHB3ZXVGGGx2buDWbSocQ8Rq/3
cnsUMoe683B79bKjMdzfVFt4ccd42fNf8us+E9+Y4Blh61wPmnQBpQ1ZYciWXNQ7
ihviKoHj9NJk6SF4I5h9GaUAO/upvFEndfQpI/TDV3gpQURTB6NbSyunqg9tS2wu
3SkLg2GGjjbPdZO+C6k1SXzXtYS/A3GpEZXiz1CmwgI/38ucYoiSryoGJoTcH9S7
Dsz9eJeUxFRS/8aZe9vexqALgfiW1KfVZpx7lxsUVm3h6I5AIWlJgFozxlyZDlYW
0fHZTVzZmm64zKW1UAXrIWyEleQWs75Bs8ZYsUtGZuJGaCLhT16vndGbGuwGNNfp
qfjEeRl7b0w/U+ffLz8VEh6KzwnyhJmn0yrXk0AfYG9+752IDQPzyfFHJI2p3aNA
rfA7N+cRdsV/oOECBBgNxQ6ik/3T6r1NphGIlZRvy0GhAm3wXY3+EiF+N6Jj0DGg
QLfU4FACap5MLlgOs46Rxz6ih0pomCgJ7KX+uRLiy7T/yNk6ks8+oBzm4c4S9SE1
XmvEtJYwSVbaXS7AozDw8mclRFZscxkZP46uQJP2keaQYfPiLWJwQ6RsIwFb6P1s
xbyNqjL2U0p46th0TpPHz/JR+B217TIX/inLtR01NAyG8sohPB8HDv9vei8GqR+9
PSAH/9Ey6i+IPcxFYUa+936IMLUlUmCatND+GunPJFiuCZEThw/sIVjCuYmZMu92
hUGN8zqMvNhsT4hsU5lykUzagOVludxIi0s0evxZBxuGMcRG6dTfgniMJEoeM86H
enMkc1ksnrBjgxgFk0kDKI08uUfrs+HeXh5DxURing2pd+NnbghnOnfrtySq4Ziw
+ebWKQRR1s6xqrq6oA/aCvEv/UjQVdIRmkie7kuFR/Y7jKI4S3cTOKA63puoCB5n
tgFXTbW9vsV2D/qRjPZpAEgFK8q4gu3VOkAcDqOdgEBciX+PD4zXP8s6Css004ry
KhVSb0+D/4LTx26+XEtrB5Hy8EpUMXVmPMe65tzvD/b1r8mV4voIkpxP/0HzI/Wg
DkLmesk4iP6aFcZ2vUDomoMtIMfNdqieKfUukAyx7C2zK06VC+G+zB+EzbttBEjn
utmBaS1RDh/oMpN6pQgqSBQUnSbCOhaONMbf193WKkN6LMIBQPiuDNS1TPisbOzD
D6H9OzRvIwx2XfqCxd1SZD0lqiipNI8Z8S/G11d42V4oq/JcKoV4jL+nyZ3R1kZg
I2vJHPGbJmnsXR8NbJnHYs061pajzv4Io/tsxRWz2mu4HMJkLs5/2MSfxf+QbfdT
PMNKWKKS3X7k+13exIWtgeRKeeLDEjBK7H6tbK7FfC0SzRImEGEQmwIdQm2iuboo
InMaZwpIVVq+qMgMXBuXntpiCHltZ+IpF/QZt+6Cu7BhljH86gUfd3fyuDkSVAdp
x/XB6bSOyjo5bE05pVq9L/x7zzsr783xXFE0meGTybTqe3DuB9KsefHq8R3SWGw2
5JAh+5HyVnrkj4+W97daNLDbaXwc+UIZRiv2to2b+rgOMfE+fJoWbkAXxA/1ca+i
Pbu6HPdjllSDF4IOlnavXtsjd+8AdHHd4yAIHzFwtWFmadtkn3afwM6S916FWLL7
jCsbKnFFrJdx0QZHX1N9gOn+1vKLuyuKA0QLtxkvkuY7BvOSidUvc17z6wYYRMfk
cW3Gb1KA61mCeoeSrwxUJOeGxtj/9FhokgOcR5flvaJy6A5hyIJwBh63b9cPUTcL
mCh9GHO++NYn4oxDLnLIM6W0fHBgsQvWpTonARA+fCY46l4KCsE8a+2pFy/pL3/j
f5EQPY5dOki+Fa4nfckkt//fPCaKd3BSKCaWjozRh5VD9aC2AXdiZbANdotARULa
zDdoYmAFotqGq4CxhCF9D+sausWoW4HlkSmI0PBg5ObYHEIBOw6cHp+DIZaSbtHz
Dml+n4geEMin2GZdMJwA5vnxbS6yKSOv5KSfPESB3kmU+7z1tiwg2VsMBzTxHrKo
jRE+4RGZHEyLn20KmTXt2WX/xk+UGFTRQxhhg64AXrgNXqmmmB6jpzLp76Jj/9J5
7GEoZfumD1FaRnQs6bu/NobLAk8KC2oaWoynQQxxgsvhGqpaRfNZIaSY2ru2ATWl
n7RGEV+tJV5umUkJzWEsgnscw52bmO8fLv3T7SEDPG1MY7IoVPtu0Ta+faw5Wkkz
b3TYiPmgAWH+I8LiVqd4yxACvIy6DOY4OeXV7qLiYBMg/nW+IjQOPT5k7Bqzmcxm
KzIiCsOwAB6IZTzY8zWGYFW5ZaTszDMqwbWqI/JCq14kVo/5IsLUCa7XIoNgleGW
cfTARkcjPnhGHfHxe9DsuxfkDnHug9XGbzXTURAFj0a4kYZW8HAFdMXYpyr6IItH
g3AGy8VUSDSALBxsXHuIqRM+XM9ww9FNG4UZetDzojnBsRgmlapWasOS80qDh7JJ
Ag5afBxV/qecPI1ZCf62FhOcVUJjbZTkCPfMunq8hBcUAz+4FZEJPjjjVFA/vsu0
n+7Ut9VODmHtJo84RQ55Vy6WWhc+7Qho8ja/exRTp2LjWuAZdMtpdM4RWP9CLU8e
jmj4Bcr9goDJeWAnqxfUp8UTw6BZZ6EohuTW+Tknbekl1YuSy1hb+RIsG9fljMnK
9hKD1btEvuSifs0szu0OEIPxGb0qauD2gh3EbJvUYHkNXyVEkNlofN7xGF1mxKdR
xAmjgwEBQgIKnegSlATRLNyBa1AlBwDj78dqe/U/HCHYrTFD7GWH8oB7tzzEzfFT
Mc6XO9H9CUmABAIK4tNqRQ2KO7bJIwiuVNl04sek7r6YkpGx13h7JZeLh6SJ/A2y
SGVPfiMrM3Bjk+l9JZ3YALoigqs7QU0jb+wQ4eQiJqdAXSRCe9UbkjT3KlMsjTl7
jMrjewpJrRicqL2qhaDCgLPsr2XezyetYHPvddNgfdUXHqccqzRtCxJSPfHRdeID
U+sIVfdcg8Bs0PzmRjQkJRoiEYMy2rF7OtnTpVaUlNL9wTgUWYvh2EEiJLuDKj+o
cSxvyzU0gtjqmbYcLkGlSgAhAWjGMU9eEwYJ85f9sfrdQPKJPTFmy/C5aPsGhyUg
I/QxihQ3wHxX9Ik/fhd6F8plfgTi5/XRKsg8HSHJDqCIito0U2fk8yS1fYd4gSmn
bmoeLy6dnH6cRx8hbaFlqa+rIVbVAtsOP3rj3fQ7KcVHl7u4W/0Ul4Yx+46x9jdj
7qmgzQjbXtOBFE5UTCCTtZCfD+aFXPtQf4PXmS/JGrJ1Tu9bR9Sf4Z6jrWGdnDFU
cyOcwd3CAbFSVmVMaF4LiNaKqiOJLb+7nxuqWWcIueWfTSYvt8HF4lcOs17uJVDl
4bDHtwpwV9QqpzWPK4pBvo8Vb/kX6tGjncVF1rsQT/FMXW5PYyXXzw6qcCsZCG0F
JzkRmmetj1H4LZPxRguT93yk7ZE/mqym8XoGa/K89vo0cdZNbqD7iswbB6U4BHxm
JctroWRCTZ9HwI1M+7/xXWFRGv6Jf0+gTGhWRDbjm0E8IEgpU9GsqGwe9hr199zu
qAuZz+FQctaSjeaXBnQgPU734GWXccYgbzRAoCpWWIA7p+kg84fRhFS+plFpmyZO
negIM8Kcr0e4Te2QuHaimz7onEFNxKLYWt78ZE2ZPs4bT7mWdHqWVrMy8uUOMF/M
eQ6MjqLWjKaaNVGqCZ5MqIox/kCuJW9F/IU4JGMCs9Go52quvvn7TAVaon6O9UXQ
PUb/XpJtTu5lDSY/uNkeh2UW3i+MhGNXTu+Fr6NgOiDf3VOmMuhVeaieExwAoA5y
WZCLneoVIjsfOqmvvyUjK0PDMD8PmbCtHjvevp9I8VrASV8g5WQ+w6kyogTqQRs7
eWtX1DuoYpjhS6dV76jJFk6FlPkiqie7sU3AX2IW6aTg8sTkNE+PoTY3G001je7j
XoLzJf/e2555WM3Xm3crzMk4hgsknhTuqaeF1quxAK4Vb+OhmGPDBD8WgA7JK0Zm
ZjjfHWTziD7BHJf4ZP1fMctnjYHcQRJdnsxfSlstYk8Zj/RKEAG4dZZb5IhzfBoa
f3byhLr7FLyKsUUp7hhZd2Ch3+mZ63krdGqRI0/5uJ+HcNRTHViyGCxVxJW+gWXN
8OPOKJ7+8E/EdbLcC+DmczlPW1lycnZz+qg9fI25MfTnIL92XtI6HQiLpGdJFWjh
aQqkQ1TcsY8b+PwvY6I3blWy80V/yfkdhlG2zJd9pN8ZamgCSt6PXlWD4JDVitV/
fWXvTGN1lHGroLeJJGkKiT0Q+Zh5drmSZcWMsyXk0qlMyjH5p5iMJ0x3TF7nlPkN
wkZ4ulkq7zJ0RDTLClixPYLojg797G636K4yvVZcxHoyMxjwjWwoe60C7dVZMhaO
uafBPdx3h7SJLzF7AOlw5pPu2LjRXdql02SNbMJKtlcnPlhyBFn2U8/ScVy8UnOe
8NgIx59B2MpKGhr0QeMDSdkOG6fhDwD7k7m4XTVx0Vh78Q/VnHKzMPXu3Vo0matb
MHTm9u3efMIDUe554/RKZfKZj3+FQMnDhJPDIQg81tLhhOaW1DSRg0OAhC0W+Ajs
KuF/1FWcx/GnIXvoM7QcQn56PTPz7BaMAXMQwse3uNAnr4aC3Bdlpdml9ASr4EGq
eknYl51Z+PMXpEG7Xp/mngnKxhM3CEQ6u8pqY1Itx41nbgyCoStJHQJGdFScJYRO
vYmNbvg7I38c9/29fUJEfTYdl2VxKtV+tTTgmPn4Pp3nt+sZ289USTtfvUamMklA
1Hs1AYAMe3OWVMZO3vSssq07jcO1p0EJjs/+d9w5VUQBK5uMpClbZqDC4++nOzN3
qbth5QlYhgIxHBdgHX82TPMTd+RUT3zJfG99NBbosBuibXi+rWkcHcC5MZaVVmdy
eRhzIB8Bzq2fCRv4ejXvDbcvwa9Cxie5nJghMrqWT95Tqi0RkONhn88PiBk+EePS
wV0US6Og/X1+TZoaz4l88q+7Q5v+b2PbM2dCmb5TtI3W8/LlKgbd5PlasYQF30Ek
XiW1VRddD6xvg3z+U4xKHpTGppadKCEUxML50ZlDNzPunScoGqyhr+f5UpMyfaHp
W+IFNRYnq/JBJhEfQKgOtkaJcHYHvjEfDaLKHpr4CsmpbuFLEgoX4FqV1R+RoZ5H
2UHeHs2z7Dyc+gBCGNxC8jbUgE0ZlFefH2sOlbKl2WmbAcESuccbkVZj2hNi3IjB
2ZKeaqfZYetw8SE8lo92p/oZKDh7M81o09OrmMkWtKIstxsm+CRn8nFwImS5Nvyk
Oeh9oFIHUZ315WYobE7PoTmEa21+RJ5GWzftywZKn5X0vcxBm83BmJiKRqQROMDc
tUPI6oxvdiQiSSoHqUSU7DAZuw214Tz0G3Qa7Jn5sKvoEpdQub8RM26EMIp1WGBB
9Ih1bHWayYNudWSgluIa2w94eTUX0LuidjFxiaeAJWvfTWI3aZdBojo0tqyUHTVC
SCQ/WSVrdh3lcw8gi/ecbztbGQ4rHu9Y3JJMRT0tfalXsYrUYRS+TibtxW2IjXQt
TQ2NXc1tFjK2FwJ8x0ZTq43tQFkM3/PP7vCjPJSRd7QSLnmlaMoiSHNyN6EtVnT3
i3v4Wsc3szSgrIaJZ/DFcIMYQWeAXRaYsIdy3/m7VHf6Q7AyA+Pkmfx22DOJK0VZ
7exgdGF2nIc2rerFNh0AAiM1zKhknXGcB+4560o44q/z2Xc+ZjFbtuE3Lig6HCMJ
c4wtB8IhxJKMz6WWkAfnuowj/IxPAwIbiUTSduuetObsyGVV0WuTHyOqinmGTV9i
BgpNXN+7Y8ePAznD+QzgiQf5ISEQnvSnHzkAFliwp7FSXainJy6lJBNi8pGKmBZT
TXcHLZyMgH95uT+1INFSq/+uwvgOmUcNYXNa96yarXxG1OOiLJsu3UMjo4082KQD
Kza8Ir3WynP0kS/jm98MCN83TJwt7CBRN539MkocW79aUjY5gM3vyS5mA/Dku2h0
Uu5XYDKZdMeQ8ql4mkr6Pd26TCoNtUV1+SziJy4bLDp/QZDogCPD9KS9Z/YEMye5
+OzTx6Q0s3IGgnnLm8qhfKhAOBX2K+AkSsSsDV+UpOZyAOjhjmTelCsCobJP50iI
unb9EUR4KKhiH6eMJizFpYwzrFtnTCkcUt2SlRXQ5d5HtJ8UCUXc9Dzct4ZDTd/c
6293XHGwK7VwqYL8suucRZ5K5CV8e1QJxzxCp8tHtnTQN2yGkg2J5Drbiu5DgsjK
3Hqq24w7xjN4oUM5LjeeAWJJHbu1Sjt+EiyLQPcdPgX8DxkacYTfXVZaFFzBNcOc
ZJ9JOcR8zo/laZt4Cxyn/AtTZrs8wjNy3K4dkkCW7WZz8k6fjZnVi2P7GbxNkomV
+9XO5VpqjcBH8sUYS+2iHUlE6g/Y3f9t5ssUhnrFfAha9ruv3oHVqR+rQTfoc3Ow
QizORTjJDm/FC6bu/yLZ3cnF0hcJL2Qu2XIMarp1avRADeNsRCm5VnzrhAf4DGVM
v0hznVc6vGOOev9Uue3iX7e9V+EP+cc2v9QG8lJLW0krEIhLvxqeqlEh6btFiJJU
G9cfsyqx4o8+2Ha4yu8X1g57ahkusTyqXxzxKBo5+urHzWCiXnF6MMM7BCwIY+Z6
ic7RMyKonvL1e6HJATaO02a759e6imqy3bkiVVjKiksIWaJr0pmJknreLO2OSm/y
w0HMhGxvuOC+V4ZJVAanDqd/pTKlfDNrGiEj4H/dExyoEcQ7+AK9OcEZLkyLddMw
qy63MmGo5eItowkM/kFq5HaLBL5XvLFdf5weTXUJNcyut84oHd1YWk8fdrerhaQF
w3S28ei0xQfYog/tUQg1m34udy46WjudaCgTFLPCHwNp4u2Xl5XlnBdO5+u4vYa4
e2tOS+Rl6pW2L3NPOqEjoPwrOjcj65MXs+LplxHL6qTOWZ0yIxIPL7y501U+FQEb
SvNfYNykSdCHauKOZqf1oku22FhhNbrdaaB8qvChQ5l702Oe39qnbiA/boxieGf/
tTLqE1k2UrOXBoSgKZsZ7zh9kw4CTPrHBg1r9Z7luPaK3y1n6wKBpbdg0VOxd2OM
BoTt2JyoN0Wjt5J6qMj4t8c7EU3n3oLv8MAhd195/EvYmaXtktSU8MKGcVWQdkIF
TlKNAAYC+p4lp+hvqi7QNPNp/MJ0pLl0ZzgRG0AxY3FEvqgD34vuy39LJH4tOlmq
PNMtWIU3CLxN5f9X2zX68eadoVxCWxKa0ZQNwoDvkWeTQeFs4rWJQFDHIaUl2liZ
rnnGLxbRUPqtuvhq15tfzuul/X9hZxhjZxymSSHdLAuU1KeJo0GegDCKbXlzX1mt
oSMbaqUAY9U58Wr2eTL88hsjgHdzMgS/WgzgpEOOGLx4k0Ek++hts+K+/xOT+91l
XmEpOFhTi9gV8ViRR6eHb6c+94V+NWD3h+DR/RMuMt6AH7/gI2hcvc8pdCh/B/jy
Z27i1cNXhxH4h5lhQg6sHyqJ2oL1WW9u+v+IeogQbsm+HAAPUIak2w+ut8W6U8Bj
33RX/iOYtWhYEaxy6oztLfMjlcKLGLFkJJ9KLOMB/eaLq+ayK5lfdBbm4vB0OJ1Y
3EiHP03qzILQw1VSqdGQgYGH+VxmA05MA+A3u756o9wW6GVtOnQ7lkReGxln5mrx
NmbSALBWzmwAFMEG0mybuihBuDOIjQr/dj+Ua/G41ivMf47EHD5g4BC7zg/h0eQL
s3L7DF55TawTLnJv6ACkznk2tk1JYRJvv8bpm8p6VbFuOeVWrPH1hqY0pWAmNZRQ
d+Z+b3BGXEaWJij/GB7LZ0Nw4NFXVGyd9/iI7iMZpppia+QRDeTfhiXaMr5puIZF
qnInLRVOxbM048XCTIFCRqap2oxAaDdftZygl0kD262KNFDxHe5n7zkZN9zHq2Li
G5DPefs2WJQcQt6mzUsaUtGG/DqGixmul4lgrrQHtplwbkO0vFock87v2cN5xm/d
tJJESIIa7QA20hSLxdZIk3njnXMCwb4YYmPqmPpikPKibPIFMjsWOaV4SEaSF5cc
d53YyK79BRYIxVyHb8wIVPGMnj9SjpFrRxD6P8nzY1a23xL4sR3jBvlDYw6tRauT
MiR/3cH43VWTuEAyDLWaCD3IOq+dP3Y43WTqUPQl8O6xUeUNgaHd0PjCKDGHy13q
g+AGaemseew9HmRXYb/WPv/2f+/rNzTwzK80PTbxG1c4mebsS5gVcIPExElN+kqV
vh7loXKs8ZEN++4IGcbaklSJ/KXBOzNnI+L5ZyPCAmY6n3UlSBLw3DEFXjc5At8R
0s828rSwA8hL0Mc/bkt4wW9bnKJInbnSYzKmjBrKcWfy/YPwVOMlBZyUF3D6nRVm
CEmGx2iCceYwr/CohSFBaN4SAhrEj7k5HaBgAopGrOQSIzJgyspULjYbxUrHSnl8
n+dyO7hxVbKHxCivL13p/lhuBUkg73h3noubBs0FnmXPBMLAS01NJ7KSXKk+s5Qu
0EYzqanr3T8pLSMm7i0PlgX1wv/78fzdg6E5KS54mS4PAkWiYwvjT3Tadp3vL4b0
fT74bfqzW7cFZuI8lRn46zyACfxET8BT+xpuVguuYLlo9LABUpRy293i4UbtYaRk
fZ+PpEXBAgM9cvD/WHkVZjXZYZvUhFSmJKN+3nZKiMjkb1jkimeWjOHM27Uvs5OZ
mTOum6yTS8/Qw6izw2iFNrEMKbnKXoq1q64+fjDkpFvg0W5SG4cPjSOgQuzZzSkm
2XrVFoDvAXbkmjjoR6Az896wLUn8flJ53nhwjuzV2oMlzyETTZ2mT8TG2Y3BRGQU
mvo4ELa9lCIjITxvRIUA1M8CvfcosOH+mSFpB5Q3Vr9CqpQ3pMtoNeF1sQJRIwaJ
7SKLWSj0DTCz9KpBz2WGgo55CrGlJwOs22tEi0Rcqlj+mW1HCO81yGupUPnLV/8C
7CHkCMQtEvkk7WA5aOAlZfdkNI0V4xhfdsmu3f78LkwokUHH00gB+knNK1BOFD2c
CGNopm3AS2xhg0OZgiS2hhALpHcI48Kr/xIAaZGKYCJV2Y7vxalPTMtQDN21q2d1
rkG7Iays76db7z/etr5v+oO5RC6HdyKLHp2Yc0U+oGYjEzJ9+nj1/HocE8vRifAA
5IZM82z+riVdc+SPfO4spApoP8BQtc5Vo3N/iAuJr/S3KXOVD3dtucRL1mBFgxuT
5R32m40gSP3zv1ij0pKR8uba4MyPkKOoaxfvxCsbYCyUIvYWSZ7bAjLsObujdUMn
c8pthMU28/1FewqiHO2jMvBhX0AzQI0g3xnDDY8+Sm0X+7xuuhhjZXvxYAngvSVh
JNp7icflPFP5GAaHrRdoeM2iYm68sWujwy6sMcUQmW7dptr84WS7SrDvQijBezeM
a20ds/VdaWa6Rp0NCyEj+jICNUrx0xgei/EvUMz+/nEclfHYUeoiOWdgYu5R4m7G
KT/RdpgjFf2KSdRzkKD2CqaGpn/sCSt3S8pRcwe5lDUmTwX4XTKK1aNJjkBrcrbJ
XN1nOWcu0w/zhYuvjE2SmciZeDnbuPJiBgB0CmsJP8rKnNdG54KAUTZS0zQYYFHG
MgVFRx2e3hTMI9HKwllh4xE5NNOTCwVn2sYzljFxZtjREfJGAXEQW5JQFRBugDjg
QIClrP1/ohcPom39GKJnH8IpVAAwoHeRnDQRRzlK2wxjnab3vSOewky05AM/f5dD
8roDYpXkMcQFdVUUG93qsQfNbTWxlufize3Jv5TvqpV5deA+UtOt627meFUqLA/c
Hwf5l8zeABBxZOJM4fzrV6L7ZLtuF01Al5xxja80bmNYAErapfMFDAGSh9oxSRJo
8beZkiKu10sbdybo/Ok3+edEDQLrqfyldNwNPv8NnG7rQMMzfG9su6BrWng8+b2P
TvDPcsvkg8xVUTun3ZbVzn3NYFuiPok3tjOY3efb+iuZN8zDraEnAhFG6MyWBrE6
GH/9wZQuf9LtxioZOuUZFgYR+u78TKNa17kURApwAG6WQQWOQgfd/vcF/3WFH3tt
4WB+111qToJUo5YJMvq5U1Di1NwO761DkWJ7VbDvZ87u2sA35iKtEignJo31SH1p
s2TqGL0wUmIYnQ7PimaIkfZO0weVUcXTeNvPqDatnQ4IKogbM91SEt0EzxiBThFI
TjKIB60geOey4yN8AfyOTf4dqXl8nrcai8t1TMv90SlhULd5neOSL73+RSBKj87Z
FwpUpNaKB2qOc/3U3HQbu9LyfeWSgvtzcFDVKojMMJzT/IaVY2g7mFW47St1R9Wv
5vRDcHhsayYZ/6iDbMsjisTAqdvjMW0kmOuUYqL5yAX2Cd9JgYYHpVwFuI+Tpb4u
nFJ5XNUiIG/PUn8G+CAieRWd8QtaltX1a50UHVraWZOuFtW6SNZdATiORVVvIckd
nbQnoqEPjhtxALLhRCqasLpyvgDw4Iaeg3VYn+ql4sF6GMlJtJnNJBM56d09GXAf
03mSXeZ2M1r2yvdxSucE3JxfpTeAN0d1z3Aolf09s7pM1L2HsFGUxPtyMaMSDc41
IxYaQPVjJquzjFlpoy/tkIbqZChqjBVcjouTua4foF0hs/kdUPBOTL+xAMcXQAc7
SiQJyAUIAaDZZ6g0po3QVXeGkKXWnc7FriQZgO+NuYw7A8PDwAAtTbjTH2J6VKRc
oEzuaCk5OHBn6pZDxna1CUmGWyLakv+KwXL5Zax6T6TVqwaajZ/7AQLmv+7cJ7dx
OxZCQIgV2DF7fQXdXPlU9bxU0Rp/dsy6q3QZrZHFWS/6dnyR+DiTRvvskmkiEmo4
/BlI62FwVORITfDk3lSZB6g9RxcsClaFl6+rRLC6YrSlmCweduQL3DujqcjUhFba
OSrRKf09z5fDBEME3+vaKiER1XKJH01UgtKby5KkV0e6fDFdkxSwwS14/JdDbnHX
rMPXdVRDSq8kVmPvGVfNLia15UvijEv4aiZ4jwehTDwDUw8wLPGC7d6FcmrfaoBs
tyEltMzyySanvTw0fz0deYb0+CMza1hG3+S4fEdgjrLaTbo0D0gWRjvSKJHb1ulB
iF4Lh/PZ3Hhie1sjt99WHC2ZDumT71sFOop4k2X6qTdW9QHKo8eFpa6K7LfbQ4to
kSe9IFHfTBUYOZggthfAVPvInTJBhRyn0wFlpvIJR5QfaTGV9wieivdJqdDpHsUy
xwuXOTcqrUEvp0UEEHN+dpINvvmoO9CacWPtebX5bPs/pKZrYQTHR6PITZ0y929M
sgXtc+xxa1ZyM63RpJzG93+mZF9cvjNJjFZBDMCp+exB/PO9rcssg9zNHKzt43O8
+2RxOfgiFMR6FWB8mQD8xwQgmKEy2VW7YkAdAM+KlRm84t/hnfJ0jhm+xogKLQhE
o1Pr4eZ/vt68a1hgCTkvdzKqJXAvF6j9prUpCikKjDibyZurjGOeKfOC0lDaGcqe
zg+agGdetY1W7UgnfCuvVgYA3oYXeKhhzylN3u2kcl8ei/hOYQvXLePJeH9n1HCI
bq/EpkSgMXWtWDT7H1QqkM/SVWzzA0zwCFPy6E4t6JnOlVBlBZk8QGzXWvfFsduF
jIFiyERuBTxh90yA7dHWqWiROUShrDUKreeRqwI7icJ28xb0tEvShkzh6iIVqQ5d
87C6K+kAb4OSMlRPnCFXPTvDyxAF69IHHPAcLiL7DnvdyzOHvQKcb433HwkeuRry
PJy1GRuAk5fpAwtULsFj1wqEl3/ZnIZM0CAl/gBk2iChf0BLUYO82JQ3xEA3kaUT
LYb8heqjSWDJcl9Xfb1LKD59Aw6tk4eebauJeKByaZ5Xu0Qk2iurWWSuxaesmXNK
dAnhdwy0Vy6ZXEY+dx1WOycrZ5VCK/TN9UqbRzImTMHH6eSlyt5QUxlYBZUwRA7G
pMA1kIlqbjZs4jPydTU27TCi19oYH8lbPKq9yBdZh0PFFpiNqldq9rT1fEuajO1S
5vbJC8Tk4SoujXWIX9Ch8guo2xrT1TloMy3kqpLfRtYRIVnpjjLCADQWwMX4ZI50
TwgamJk3B+d7j7sANJczmTSQtZTe6fFqE5shHUF4si0QqKW/m8IcoOC1QTi2f48o
IelC0dY8lSIG0PxLRXJbmUmtlX/siOzddE25S2YWRTZm9YBYoFiR6bzqJXDlcJpa
RDNTg0TDqL1ICb6HMnPtUP24mdEpq9I16NL/Hc0Q5TTVvJ9l3d2sS8uMqHKoUxlX
kYaqMDUUMvYcf2HD9Z2bMRmU7BgEOvswC8vojReRCI5jbrhRpt65Wdh7HwQ2q4TD
GIhhtiJ/ZA5bb8Qg73amiJfi6rNABG4WketAnY5y98lEjkkRXUUsXGp5OtXqk400
voX7SJqcGr6lrt+UWKZPi/3rqhZHh9HqI5sQpeHRG1xzOFWjMeNx+fasWz8ZTBIq
7PBA8uXwS9HqJoDlnoNOlTxySmkkhntuygyN1xkBChxqYdt08Mtx6cG99Hhb1sdH
sFkoadCYGrk9YA3WDSM+sPTlR7uTcSQjoW7gGhk99WgQRJsZoKbMOrllNKadnHue
rQ5tAqZ1XOz9MVTgVSJX8TLrXkupdvIlLaeQlcl8862LgY2uleIZz52pbH/JerRx
Z90GYiRkR1i09qPbqCzC3lYPGCHFfwRP8luR2UI7/XjhHIqRxDiYw/0eQgWy9fJx
5G2THD7AizDpOXeGosUVoeNpqVXBcc8/mNtOiDp+VssDFHnVrF4yWDi6L/oWhglY
QVZkf77+O4dqFN6lXvO4xNyXEbKoeoWXswfaIuK1JqD121dEe3FhXtWg98yCkznE
QMwLJgRcRpz+CecLv6TmdsYox45XdOCKBW1KMaAJGq1NHSULTJwoe0jUL6oTZJfu
LbclXsSkYwEscht6IuiJzf3sIQPCF6V3uFP3WFMZU0SLlcs0iqUqHfECHbBHKYPv
hYBwiCSUkDLnEvQf+qNlXSYHIAPK0fTMb0Wjfc0T9UmpF5h0douNGnJbnZRc6mQa
dp+igNs83edMg8meBInE/bH+e+MnP5GledqZOWEoIfrk6aTXoGXsJI2Eug9ank/N
hduOiL1wO9tlz3dsFSp2CDopSkIwE2ChxkeOwkREra1PtTv18j8HAkjpoPyXYRqV
Za9vesXMc4X4oHm4gfLsSjUOMA7Iupm6X0FfTsv1fWwNYtcSbclv73Y2tnOspwWW
2BNX9WehrDYXNjg8kakf4CygVK0trtzYzjeXB6EWXToOKKtJm/VPSmAK++fKMJvm
2x9VRRKtzFO6xhm/q48x1cfLGdXRKcAeI7zZ86N0BKAwqX+Do6ywnqXcWvVJai3p
TJ6PmcOvVN554vmnLGqFu9HNaB/CC8CrB5gtvnQBxIY/CktzXiTZe/j2tP8b1P58
TnjgYc8ig4eiJXLa8CKicb6y6DUXorkW7Sc9wnnQgP+ralG5QwEt5c9ct81YstiA
WtTksqYjRKsI0yuROnGwmT6iaMXrlnr7XbmdBYF6J71yoPmb5bTfNWISJGtaV06H
N2KQXQ8LDZB4NeJP01U95JghegofcesCotIare+5OJ0/7ptcSeHHLCiVsgUZ6uFt
Vc17Izd3mATOuRXQWaauQniSn/jZuMD5sokgEtXe3rwcMhW8FFGhqiTwg2MN788I
2MbHv7rXlnJVQOrKAmHGh/AKLb842PB/rr2xplDZUgULWWw9oPTEB2WyCkHXjJG7
FETltRkvv+yqfteYlN94UbWKaA4vat+YFK6K4pPNeZkDti4HYqOJSkEiUBfF2VvG
dbYqYPBO8t9jUtKYcfJ2UQFxnQpiuIJKpXl3PmPTec9WvmsmALdG9zZHV3+0UMQx
`pragma protect end_protected
