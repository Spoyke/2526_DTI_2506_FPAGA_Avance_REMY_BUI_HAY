`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UZBhdDlN5Ufck8E14VK10ve8GSRUA8l7lkdN8KZtfNWmyEnqrxMJZZxEf2fTJJtT
bC9WfzMpj8m+zzGteRDqhlJW8g3aI5m46sxo9tGjaaZmfM4SHfNeO1+UYf0qXN9h
J/WU2sAR4LUiQn29EM83Zn1PFkfaejFP4iV2TkJDRJo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14768)
2cRSefOx7AXamtuPPeYEGncfeIHx2QRCpizYJltafHQDQe34ZWXCMMbuGzl/Ku/d
d9gCxSf2keigi65uC2rW5c4tYZiQtIl27wL6WiGnckxBmeZwtMg7+ieLtkNSzatz
qQ11YbKdXv0XLkqHzC9Bo9MdX/64sXWUKX/apIEKo8sGYTC9iIsj+bMFIO2xGQXC
jkbpANHXDl1YQSeSpW7BmXqwfaNSbi966LVT+WE/aHBH12x2qWOkpXSjbZZ6fjl+
c2UjbFF+00/ML5bpZArkVlM+gdkEiKZBSW/xtUVvaZGCcqMa7g6XbDRAbSYNBbQm
ksC13uriKIKi4Y9UAFR2H9if2dJ0rr76RmZUDh+DFtS6fA4zgnKKX/XDZsdE92lK
PzR+oky10i0/FtMMYWPkBZTFi6a8J6feo7GbfycgNC7YteoNtXmyD7Tuxdv/6HLp
FTesdfikUHgdOx/fv+F89MvzcfFEwJcHtUc6MHeWpzbf3mwickmfvApQ44WMZi3C
ugBJ7gyeENi1SpwwDnyHzkzhxj72tq0Jl16EPe7HfsVp+dlb2OSwMTAtyLnOjN8c
OzvRpBcmefD+KeuWr5rQy9onmPMxqZrUoqW31v+gqj1s6Ec5+7Fs1gU3DcoRedIL
TUdutcLOAAnyxuNtqwIbLPjxzSvFxXHlmTHYbZNrMQ+V/8bBl1BG7GsG0oP8cFd8
hxixL77xAUTH+LtMdbIgwPQgMM1lFWG/QhK4lbnALZcInu7X3J1QazaxnrbWDguE
C04XmuxTIDqhGvcWXryFisff0CGRzUuHneO8Qj9zi36s3GekWmDSWvZBNjBL4D/H
fRwMxp3PubLw164JnoGsqAvVb8+XozK4zo28/jG3893Gttf0+nQdbGiGnBmvUtyE
2mW+w3U3IFkLCyZCpWFSa86YfcDGj2cepxWffdQj0nSzV922ZwigwQ1mQSsojNc+
KErOjjX0Pj3qOCM641XS1ettwG5AnNy9zBM0uGcI70SUPx8UGglZpNjdk62FuEOn
sPZB/XljXZmtz6zP+xAABr2JU9R3dutcXvijJ0yZiyHX06vG+WnLAOXR7rBng8VS
ZS174fO+g23UvN1ntRiECcIoOQSKGE0BGQvlCrJN8EDmpBmrbqmMeeTF25Qg5FRn
c9D3vx6h7zcRihBu6wctlDa7pTRAkdKCdm3sN/dDYtDYG+t4d4b/y2m+RrWs8gY6
7Gxt5ICv7/9DqrBilzGTpmm4zfhy3FyYNsf6jbRTGe11zxB1bTWoIn+v1T/OMKYk
Mnu1GLBTtPoFvEocrAzvh3dyEG1F6kYUUzjqU0d8A5pdg9FpRebxCIb9kLakB++a
BHCHwg65mAq8xC5k3k39kgPQi8rpfTtfH68L4y0fm+b6Q2E0/XE0l5iTOGNd729X
HnW19LVNH2m5uMBDiK0USrphiYbCKKLuQl/Oyww4WWrOn1ce4efAN54wQTjILP1W
Bn4hTHrQUiUvEA/mwlbddRMBBOYjsmf3wVs/pJDmN45VctY8sfQPy7/JSPrcfr8I
tJzpI4LS2NZde8yX5m1gDJAxfxcemDKieHLaMSMMH/2HvD/rG3Rm1hz8Utm6ashT
q4WcdZuQE9Ty3ehoRePlaU9Smiltj+O/ut+6vptbekbJGZ9mpnKLV7yPI5kz26xK
3sciXwEBHNYem4i2U9pAnPDQ0AsQa6Oslh/p4Nr4Nf08+BeXWVP+P9hXj/NzlrZS
ojwoZkE/H1kj8FTFA/gYuulmToE49y9Tf/6Dn5vyWM3+LQrEBpAqLeNcLq1uosFi
0Z/rpG3Ixm2E9IcnGhVdeirjGg6NTPSqDgdvpkNT+ygu/pEj0owu0MmzyEh73K9H
X0U69lmMXd5v6b4OkpN9IReGb0rlrRq1dx0PS4awM2aOGAfDMD56+j7z+xg/P/UO
o5bAl80n+mLrJ9Uz69IS7WSa1ThU7Fu1/UMKG9GG7EvRd6/S9xNHTa0ua8iWgy5r
2MKtzensRNVXBZibXwynSImMAa+2Tvzbbe87kG1KM1K26iSL2QMll6fqildko3+U
C2XrCFoQtd7HZUtmsilw6LlybrXw5Z0vQ802usYmNinNVcFQyXVDjDMNyLsrD6j4
zFyNKzC3f1sVF8OaZtj7PKWkhuiqMGeftWK2WWgqBIbJSlE8MoCCFOVHnmHVV7Zo
fWQy16sggwfCqbnZinfqeTLTlKiZWzPiWbhigFEANLkqQRMA0xnSyZ3oxg/UtMIC
npL/LzlCcEae6xUXDaBnbFJOc+LTqn540lfMcVd7nK5O6SxFaMKJYzb4AW6ZNsJL
VU/BhD1XBiZIvL/G6oGt1aaQGnYcdKzJhV0Wap7X6UGPTXtPy7ep2AfQVAwn57Gf
Ehw8EnUCM+a8Zyx9eaUnmZK/icCjc73TambOXwy7ETDZDhvrlDaYhAoouzXtYIpJ
cvj20w0JcygN6zi8VeYP1RJ63bRoCNzy3VIdMYh42r099fjg/PPtvGZFO7lJJq+i
YQoCJr6D9ERrow/xM2OYmtYMTE3QafeJiB7cesLgv5UcEJvAydLJdzv3WMZ6dSag
2OF0sOSJcoUfBkRBBYrm32hHMF1X17J8FfPHrl754/03vXPxqmfEBe4Fu0lTBcMy
6/BXFEs4dohQZfkHJiypaqr1v4AUR8GzdfJSqvsL5wJgG45EkBRmX0w5LNVTaQou
KqdNIY9LtSNmjn7iIns/gurwz1HNTq9J+gJx5isfmsRoqdREtOub/V1g9VazBstV
+dq4iVXlhgAsimGk52JpilwQinaiGi+eavr8Q7elHP64XB5v0M6Sz34OX/ZoTe4x
PIHA4FznRaYZHD02wU8xqquWfy7tQwe/vA17DAhPhbBytBePynguUcVDkBZhKQBD
rubDahi7z4wqSvDe4nylroeSnOYZ3m46Crcy5ktJ8JbmgQttYNSs2XC+Z+ZE5O3K
JJhPHg/n3kKCPnjkngyu2Gsg2xCEkaGKnaK2lBV6BFFjrR5kcr9+egY17ALKeu6C
ZZ7eDAU55482Rg4h+Hc+i4x9SSuuxLMi6OypVD4ac7AKm+vHLWIunAwpOcD5+DaI
w+sBLK2k6HqSTLeDbVOsfQPTfc9ujxdJip9KzEPgR4C8AZacUQfG1oWJS0LEMXAi
NMPieO+dxykFAZcooEMLqljEKA/l/bbFmCm5IIHQIEhbfCGE5F0hthJOCDR7OSDr
BNm0UHt8aRL4etn0EBI9ICBV6TaDpZcjeppploFoIfTxfgOuTgdphSMYxEJ3u5kX
0k9pReBYG8UV2xXO07J9E4MZnVJJ6b91aT88E4U73PWZ5vFpWrlWjkvuOVoO/eJM
NwTAThv071G7i6cFEClz9TxwjM5b+IPuLl22VBpq4AyCjlvg+vZNZe6ClJtGPeGf
19fEJbhNScHkFBRX2LJRydEj864CyA+dpWDzh67D1q7QsTBi/Px8qLOlckRn21Q/
m2AioOOTRfYzNysChDF2pW8IFmWzn9wcRDLoiFI8fOye4H+hEoAFOMyFYTvaazub
6yGv0v9yloOPuEMsvRw9rjrTZeANnVuCdcFUlk0VaVW+x0Kl+TK9O5jT0FVEfrGs
DnrIZjSTArtn9b0A/xm6IcgMUZUMtQaXbRtV1meMvnx4fmOBgay84+jyRXdO22IA
E8ov6yVVJiyrtQM6dCnWeD7B+Jzar1kxDMmasxYt6SUUB0X34wRJbXxQ2HCFzMXg
jYnFtuNe9qVTJDCS59j9CrtmXCLCg77qLXkblWH5oBicb1f1ISEfJM3MwmVAx7nq
vahriIMOXTemaCgP24jHHPRECCShv+r4Y/hIpEZLLHMXXyIajIeM1Yt2+5tiiqt4
kPnTUv66vS9svbi2F/rh5RjPGOr6kI1TcVksEClXrqOIInFaIV6VlLFSTKR03oO/
qQVIlqzysSwz+hwFhQwiY6whR756TK0dOWnNnpT9CZg/0eAy2UhcUDog1Ym6It5d
tvkCxoO65fqgK0DOUYe59hUIbR76Nra5bj1H758kwB7HJ7Mqdobmg9sTGuRjoPST
i5EzbUsGItuuhEADn/TxUaCj3It7+HO52bMSNtN3rTLaukeU77k1q2msi+UqmvHx
i9fU16XrcWWIn3qD7hgj1JCJb/2U24OUGBGSwuVik3qsTAgJ6CQdSPJ1EEaUI2Td
72juQFZo0osabLsyGDiyXyFYPuGVpfuZ1Da27vBXsUZZSbyNbUKuVI6phSBfndAi
ncx2xpc/EikJqGjKz2BiXSL61eoUnC8Ao5+xHG8SHEJuj2hsbr5O1WaTaUiaueCm
8NAnxZ+xbiAQKllSXamD+RZ8U+pCP3agrxG4vwKMGzHUwe1q3hyjPldKSy1F6GhV
ra7xmHXBtfX+vvs6qbHne05El1jSVhnkIagtJRjEv6ghkN9o5Esb7rHqvo/98CRj
2c0J6QOTsHe2bsY00C1Rs3OfncP+Dre3tFhcAZ2hXdb1NR01X4Rodr64LdXU2F/U
pjxWpH9J48va7jUDT1cFR5TYHjUf0X9uW2Atv17DY1JS6j4CDxTet3d6iU7Szkv7
ymQMazgXF4fZGXg1yHPsiwjO1N4wEyMD4h9F1R1vTyHPdx78tNxNRmg9v4gS7Fba
AYuHDHOAdGEbsTJBEi1hoxrlFc7IMaDJEGqpuCVcGa2GErFe/2bHWkr71F2wJzJS
glfJaDQ4nFpM8jRMz/eiFD7048+f1tDAKnfs2ZFijp9RymqyDfc3CC+p0QWWxyhK
wIb4ocCFHF0dvC7TPcF1WU8/cBWA+xR3qH5jZ5LpCtyglzz8kzR8NBoR5UR6At3Z
VyjZ1UCkT/Zbfh0FcADTb1rRl7anYngFh0EgrOhRgsUkymh2qB0iLXkvooFeSWto
aQzkitGWF8Pm6Lyotf6TbEU9qTR7KY1qYlSv7ZntJpIu+TQSqlEmbgYo0f8rRIPj
61MSIGa0PFTxE82bBeo0TOMej+fbgGEniaI3HIMV7qXoMxSUKjTpJJfg73m/5Anu
YGBvCafchjk8qB6ThY4a64ekIPbdeLNB+b2GylA6ZsOCFC4dUsvusOr/5BjEQVhg
8C/RQX6ABnrd+Ektq+NjPGzUumePM611Aog0uP6bqm5rvMejp5uVoXEDtVi7MXCB
3Xiey3lz7PamR7e/HTSgysRwzICe3wFPD3aTcZ0TZpW7Rd1vcFx5e9CLIH6Istyw
KTQu8JYABkAWJ4CGy52TqqHiSGqV7nBR606vjJGv0VqRpcVPrAEP+5JY5aw3GuDF
yqhmigU/jdU5B43gFMJyQqRktJYDS80FW2CQHPD0VOAtRImQ30ICdTbMthXdXa4u
399kFqnEtw4xYKfmfZ8eYMgZQqiLKS7dFNogMP4XARAkSkIO9J9QWodv8eB5JX+0
ppBtoRGmvDnbqxIa3f9FU5CiRBtXXx3OiZwiI9IcKmS+JpeUUu1MkW0m0WiytG5H
TCB6XmPMP47iZn1ZTSmsHp8oQVgSAE6xxt97ufP5RYKdaQ15AOfwIDdP8TZCrbaE
t8fsPqHHwa0To4n6PbwryVr6yfeq9UNECAtU8Em+h3yXXoF19eZLzPP/qYNU4CYJ
5M/26ibIz3hXRE8h9DnGSEFsCKt2pNBDBtulXSttdoiF4JcXv/MMXfTUwMxd1c6s
h8dsRiPag4dLpPsXTyZuY7eiCvwbK9wi2HEaw99kL1elmzWhAwjc3ddAzXpsdG2D
n6C2gRalBAkI/Bettki0/4UjU91dvNYyutMLJKzkoCtE2IZClUgcZ9TRuguRzOSL
Qmr52qhFp1CoEM7yLzWxrx8HkwbH1WOY/j660F9YHEP3SgwBmOmw2rK4DnWXXv/E
P0T/21iRumLOGOcuFBr1rO1wjY1uPGXnESXj9SDfm8u6AdjLUluUXZEJTGw8HUc1
940montTYseoY9mGijnwl8OQMFnTPnC+xOmjeBU3+G6CyZADRa6geWBBB6wGb9NR
Q5gupg2nFHE4CeJq0N2eMfumRdVqNVwNsXQbPBe2TbPO+whvTYd5sP6PGk+4yc2n
t41EMW/hy8/xQhTZufE066e5hpJhtJQtp7ZCAsVFkwS6bouVXhFcgjUI9i90PK4L
h5n9ZI5mPyJpAhZaN2gH17X/5Mi86hZGd9iUtm9xN0sX+aZ0yTb3AUuft6k4aOqn
gimEwBPbH+QRJ6CMNXlU7tuktyoyzajSlNLzmFqa5qOZyLM1cNK1PZ7FgWo73IM1
ddv0MSy0DhC6L167AdEyoqdJs52UGs6Q++3yFixqLNf3RDPULMYoBxZ7oql5O2An
sp/5v3J3jBpnG20tz9WFXAyAbSsw/BPMVuZ9FAcu+A5e8V5MbcEP1d0r83kUT9co
rP2vfuGhu0hoYmTeRWzZaLYesyWBbN6m+ynDbZTntSzABTWebtUA/8prNAhUX0db
EzFwgPtdwzCZkYcYnQTOf69iHybdqTsJd/YeHQzDpXP4aAuYJVoZ1vnroX1v9wE/
K4nfrgqrvSfu5fUyLBuJjTDF6TQTXQQ7JNeHZxO1LWX0woaW8HGQclcnqlucQyJF
Dp2NtDKTJIDjEwNA6ozZ0+GJMDwNAK55p+mzGbE29J4z3x8IchN+juyxx79wwJi6
b+MvS4bikPIhnn8KfEuF8t2ZbJqnH81cGB477FMgFd+ZvFLMUiPIlaEXhl/1Il3z
BNLO9gROffgq954u1eRkYPbcgeWDwUO+VxIGgF+VY8a0PvJhJOVJoTDQ18rcB4jw
1lKnydvJz1PUq3ZZoq6aseDI9F+XS3FyHj+bVIuEQFrp4E4jnV/t/EFq7tUjNFwJ
XB1Chrr0XTA36l/d6TZNW/2K9xleYRyL895l0lGceWduR+SX90wPWPA8UbYQiznG
tUGP24XOUTCjvCupGi02PGHdpmjQPahKcevdxfPsylZlqw7ZKHcG+XwjR57fg9d2
p58vby9QbCptQygA4Ek5ok/pB5hSIMwN+Gk3UK4qnOts26wXB4lLV9/hR6a2DH+X
xVbiljAN3OCkHd3CUJA5BWxh2v7dFI3a5ezZHuhIRe5Yy57UQZ5Ni+cSGrw+U6Gy
IxXd7ZRMvCjkciYL/xclS+ZjAcWSnFf/9Y9DPJtV6cDJVL72gCJRinuRRCQ8pSGG
mnqydELU87Dq9uBzJwHwQaSIrs2etPsgc7qFKE9WN1po0qVVt741mjjZ6V0ywBIo
Rk2+Q4ctR2E4MswjdTB9Ed4412ybsP9XUxCWhpin2qLWdTZROfgVTgR5o/lZcPwB
fQTWTOIbZK5QjhGpcd4lGdweBnYLnYRF5TfOIVJemOgk+aOc2ulDRDRLrB7oiLfZ
nAVyX4LQCXtYJVeGsFt1yapo/GCzt1SSNsp3knyYQBCKV+FNhoMhGAu2kgf7jyFX
C6ot5PCPbcfwWaYNq4RgdIKefoiBM+sEjxnHzLtgCKhMJQ1wbfxGsmRLtcgdOIyA
wvh7zB6atiS6NOCCtxdwr3nGmYGFs9wgFZrG9GoO1uxBa5ATUlHj0uRGmVZTv99q
SfPOUT9YsRI8C4/ubSr0EGGFFsTNaGVBIePI00Nz0zFB9l26+icJbcD/vbyceeK1
aJ/nIG5qfABivKFX4zH51NUJtaSCcI1ohNYhiM9zUlEjeneDsrEJexSGCwnm8oWh
dV8rkvLJM6cV8Zu8nFrdy3JCetNimISvLOVx5fQs1MmCyjJlA8QfOV+2CUolUA+h
hmg/MdrTOhcfuKXdVaMxKzvpOxxBsx6HbVKpwIcfn7dKXUwbvfuolMkFz2NyE+/u
lqSUgpGv/tqQYEo+771LpiLHp7M78XUop857y9B3RTAkfasavVfNI+5sUP9XVQ2b
Kkvy9H2sSEtolfbR6XQOsRKoTiI9Iz1jKOS5zcEyQbUyr5/+hTHFJswv0HzAxQ2B
8uYBeaSB7vuH8e26gylgwQ0qYD1keJ9j+WvgynEHQ9JpJR07dVHj46LMBuUAmpL1
5B+n/coxTrai1lgNvg6HK9IlocG2FrLsYuBgfxvLaFOw24p22Y7YFwf6TDApWMI1
dFplNLazTKN7pFcwJN2XkZ09Clvc4heiNJhDivdUpeXJnoaMdXwpAcvEGKgUQt9P
sVKBUULHkhggaQ7GmOUrIznzuAptA5lJ1CIOahmaQrZVjQzjZWovTj8LBFMI9jFX
+Z8MdfiTwCcWf4PakpVLBxXhtg+bbXx1hfD2YJTbjL7EKDMMMVTm681mCQzOdM52
+4bzZqewrQOnBzWxvRQ6+3NXzdZ5rYOXR+VIIPBv+MmeUkGJ+5D4fZlSZ+tOPiuP
775Vcfj4IzVSleXUv4CjW0ZgXUGH2Tlo8ehaM7XxODWz9p9SyvGqou8RO+/tvCYu
aUweZ0gTcZku8QfG257OUAlRp9V5y/6WrsROTZZiYvHT/7Xw5jW6Sx78kmX4GEpi
OHKv6fnJ9yAsyLNdLv4bJxRU56gcXwGusv9JRbXminm70CBnm2+zR5RuH/o+VdjH
e6GaDNqSQ7RB95L+nO1uzF4lBjun9ZrLbhDQ+GmD+Ph4sWR8wsE2MPSEENZc2Brd
hz2mZ3KlcJk9NeYwXeUwsDhgGuzOMXnvBrwW9O7XqU4H8fof6UdrTyvUczpPAw5a
/WnJ7UFyGNhcuEq67PZv0CC81mddK59GS0lAjdeMCJdKRSjkAcKA1Ic2MUv9Xwia
rpe5Eeqb8YI1/0ihMzJrjf4m7ipV8kI4l+tbZFKMglnVkyiJjkyljoeQ59a2DItN
FkwS8OVGHFhhq7uQReCwYEqZPf53at/zHNu406WFLeccudi0/g9ZE8vsxGvf7+r/
uTgN5IPO705nY2bvv6PGpf8tHYvMNZzh3LhHMdSsUaVg6Gy1WHbQWH5ud5VoLMaU
mLivyYqSjFlKNb+n1S+MHs4IdLn9zQDOqGUI1Jp/Rwyt6Fu9IkytU6PIgoopmPXl
25fU/PFn790avuvTmK0z6b2jQOlRXwhrg+48vKM9GkjNiTKL0VuqIZRJgr5uigPX
BrC8ymC1t6U1TUbUWHggM0r9+cxtgpNa3/MefFtxHvg1hS5mXo2S+WBgsf1n4baE
n/m4xZCn4vqDUKJ59WaCchFJf8nhSAGxw9jg/AmzQgt6ClL7VsjII+zFAY+NQlZN
SQzcZ9lrRJC7uU/r4L5ERxN3z+Yt1W6VDYgZubWTkQhqh6PjmrGXzTedp+xj711b
D3SYk88ZWrf3cCXPHMeDlzLgYbICX/BjeptOy770vWTGCb8aX0cGBOfpQP4JulQK
MT40aHf9132oxDkwJy02mCzJ0PYydCH8EoqNh7Y+cQvypL2SFYFoRPUgPGIdl8CL
1w4eirqGcFMviODslO9DZNBbS5NhdbG4FHVS42J8ckN069LcTEOKnTgszSm7BKwF
FI4qCsIAEJkx/fnArAaPtQFcrYr/iTSuIt6HEQKs2If39lm9lQyXoD67mNLt/thc
ydmnv82GQ3eypfiXgtYZ5dNb53KlPqUuaNV1t5qAkYuFmzv4uQ90DjOsUq/Mb6QR
lYONcOHsDp+TSs3kkdVGYyFE6hnW5KZry3g6XfJoqoSwx2yJ47LD0POV5IThxV+/
VWCj8Nrc4sk7WTB7Oh2Hi6OutZlCTjX/ZC1xcpwn8VNoRr8aIM5+eiJm0eIPNlo4
zKUEqyNw/MpSsvrmP9xYMPXcLH5XcYko2rwbdbyFPi30CgFxj1ILOnsEHvgs2z5f
JkKODXrf7aju7cz+8oN64raIK/RpUWoh7vgF8fXfL/D8N6hwvydQ2eyTbr0RhYiY
5gz/WX0PdowbiL+Tfeg663fC/Yp9TNXW4mAxwO31mxWeMwDzF71Lcfrl2SV9TPOt
Sr/hFXplp2lbSlxG3VmADXSCdEbMAJUx1hhPfCMND3W3x2KWtPFkfxVtsppqLQ8+
Gq9qSqSHzAQ9Bwwbv6lna0vhczLnspB73tUnXxh63fA5z1QObY4/G8zjkefPW9H6
UZLmzg2IsDvVN9pRMA5AjRLa8H/JaL4H8gedJ0DJvY6sQ5c8fE/fbOrGshIwIsk7
8l43k36QX8b3HVSYCds9d1763q2QpWjuLlfbOaetRWw3KwKuoPk+IGepcaKKlSlu
/UbvvWFx1bntKABk8zeO6OuyFUL7xZhUsV3h4KZz/OLnBuOUHcv1JdTlS81uTl4Z
y3Lu1MBDci3mUtaXMW/33ZU4ZvlvVXNqB4xVBaFOp6vQqB1E2kfhEa7Msaxwoxxj
JzXbzAAq9U93FwYTP5sC5p6aKgLApynkuiFFm7j7VriINqH/mIEbfRhERwln6Jle
qEd1IsuqSGhF4XwnB2a5DDDl8AG4Ohgfk70y6tBZDT0qytcVdtvjaALsBIzhDy0e
Ic0ugqYdLodrVO0zj00Vy9ZtRvTD5x2so2aLML5cdk6/HoY+SHIONm2j79ryivWa
XVhyzGUFyqoZpr3AlEFaQi3iuytZWJro4IEEl1Ne1wvlxfiC7kGIgg43k8BcmX+S
PoIdChmtjUVR2QDp+6iN2MrEkk0r31Y7THd3hIMgTHZdxCYUqzKgc8QEvLWKagF/
1fL9tcOSD9oWBSpQOXPrITnuHDD1uzV5B632k4J2iepzCpthiRAitYuNCO6pCLaz
uWMl2J3GrNEd5CoBrtU04Xk1Yy71ChFHXDp/mDfcCthRWhpVvcU38RjN9FHAwH7a
gE9NRCaMXa88T9N4QJh6oG5w0JkS0HXNHNoCXysyIGkW87NPwQ1/HkQ1QWVJrFgx
upkC7UjMOJcb+W1j2j005MYFKLCDhpvUaQJwykZKbQGwdbbbxCplu4MlxXwyJ/ol
pmPVB/SC3eHrWvxGqmKhsFuofGXjNGKdkTXp+7AMl8mFCOPLgx/9rtciASpSJvw8
obag5aMo9/U52kPNp53hlmShb1kk4Og9uCOZC3/DQDThk/JpSeeLkbMt7m5FR+Ng
ppzbpd9qj4dr3+EyWKbDk6BCTM8DzPFAmghs3+mtg4w2tc0Nj9rkSg+Y2ntVNc0U
YlJfaZHEOoKUAMWRnAPSH6klPYlDZLqF3HKb1LwejXYku+ftBdsjzp/Oq+tXHcqy
lCCkGkoTqdI/BWvGY5lVveND2dUCrsDiRQsWj8GG7bg0TFwfFM3D6sP7Rpt0yGt0
qcnSAZ19EerZehqLBK3lhye8E3R0czcta+Z4UgEF5jhtpGhmZy6mQnEbVIAg4gSd
N5biTCfVJ4BARKdJkbayqKpE1ApNMuq6svIBrEC5V2nlgt4zlJTkUAyn0qvjPVHe
w4gjMOY3aYJGFRfPd7vQqSugeJKeFpZUslFLI4wCvc6QC1zbGpQenakJvcc47aii
calFiwEP3tcpLpp4uPhCVpi7hhT6BHbjkJBfl9Tdxt61EQ/sxg7NpAJkmBbwzCKm
F5PJEHLoFpSyuEStjnD8RcopC6qf9AeB0Z7EAoIkLwe6H6qQd/IjVB62FDHdU2xh
bxZ1TySqN8+sN+sAc6A3N/B+6kKTMlQBEAclfAp0DuZaCtWA7IXwx/DvX8qpyukC
/ksWnKpxQI5fVsJh01hE05wJZPmSUML6j5wL5tuhGKVrFJbs4ZocKECV4pGzhiKA
AG4oCwWL8LwlXBp/PCi9NdMsFF07jLrchzGlnABn14mY8bZ9KW2eiyshngQ5QTOM
UE0nAnkWf9DHFOOgc9FyJM9diHs17XDxFxnRt30kgBoOkv2SGxH43T6cuw/uBxyy
+tyleB+pj2hfSzbAomv4cpEAYr4N336xRo5T9gvja+/dqeqqeF1mfBj1LwDj46nm
GiJQQwMBe1erZOGGRrsj6S8s9MhdXMm5YDF8VEiFW7hnR8l9RcA1tw3fP1RODtjj
3nulGCSOWWJ9SsLryUBncoMSUuagMp5Ry4wYhFLBSJ+NDx0PnEmTUJdZYYP6vwys
r8OrtvS0v4VQaenrrRX52sC6ft/5Mn+HwV+ILxfQ9J4cA1vtEtOLtzoIfwxjsgEc
IwIvD628v7G7GpiFhestzoJZaLuJjrVscErV7CPVavujCWTx7XXcTHmCL+lVKjul
LsSkSzy8kqVGvewLI1FEW+kNTR6YTbdOJKl4IKGh44ObZsv8o18xjsj/zZY1o8zD
5vbb+TgErrSRyisxNA0swabqm33bLEexc3sUxMSB4zCDWQM3W2kKTTK0ijupdhnP
mp4hsnL3AOHfuVkFTfUqqNWdyN10mOgoJW+U6Ni9otjy5NtVUVwFJNflpniE7hTx
atnz+c3CLRrUdGn4z/SxnBRToSBEEzyqUu2pA4Ti5hvj7Ei0YBg+WlJdrgHzSUi6
H0fWDP+s7BdFBbSireITRLCZRnRGibKUAMdJOxkcpQIXipXrCPmZTh6L/k6AM3L0
qk//ArL18hkmHbagdLOkiOnAIjQ89ydIKtJKWW5tODqO9yQv1KcU/pXlw5QTLX6D
eXGkgNOE0cZCMrWWx3w6I+AdUvuT1T7pEz6OUyKC78efcbqp+z9DWEnlZabJvzMG
Qku4nnyIDcV9fsK0K2xzjMnDNvBYwDRI8uXmzNz4kdsmOyx1xDWqhvdKePhTHLDy
uqzRQWlXvpgFWSmlOZLNr5BqqeBu6u8XgpPnVJPb89Xum2D+EKbTAaDccoE288qQ
0CyibniQZCHIMT0vonlbLGW4Cgif5DPdpjDlusB/LaITf4STJn74No44jDLtc0xU
KcDUnl5am+acN2+Qb3obh4Nkzmw8wBfvDQTVqBq0tdHaHOQNojq5hTXKwykJaoMn
9WjbR6zwCfUKU9EVkP8d2BfKzMt51Xt9UIoVbJax6fAeNTBPovvPjD8gWSaoUNYD
FxneLzQTKMieA/cY7ZWnPAGwIW6K34MeXubIim98uXwJ4I9Db/p4lokr/A9kxkdq
nvBkVelF7FR65cqToNdlIbdaI0dLwKoRJHfWhzP3awYY5U0hNyT+97kqLeagRWYa
h8Q8gVqGOOsGS0/CUlJE1mK3EiJn4uadQ9T65WZ9VQmtCo6bmA1ABeDySIkkkeqs
g6sV5Me1nlHRnsfGoisZj1xlC/aLrumYHU4vMHMSEQBEsP+4zx3hs46Wjb/OyMoU
KTOJoFWrcxKD/y+c/l0dVVlhn2WZjiMLNB0jVaaqos+s6bCl+qWGoDQpgdk9u7ZV
fHUF9rXMEI3IXyephUd/GAYzXKjlufkr3W0U9b3O+SaY9QUfgXxAPkJCansel3Iy
EyAc/1LDOMqY3xjuvKNbWLaT/K1hr+csq2zHVuaRvxsYD0cDA7CqcXjc98apCMUA
9Tgo0GkGZOEvEPGR5ED6SGvqBnLx3PtdhbWFv6/nQXICsdV8y0DlpM16hna43A3g
x463hoGrw5TpoDfmHOQkoB20ceIt5x6WSnx8kziz53yVfzGIKnWArE6P8QpQ0GZj
JyWuJm3t68LrVGSt6LYmKAZJ282m9QTM3W5uouP6iFxBFFjSG90ovXdHYC9Ss2Bd
mA8DPLKERhiNsoO5BeWRLSYON3AKvoZAOobOOXQNbvWv6hGTHzBr4oiuV38dlbY7
tn/jcGEGF0eYTXJsJo8dORE+IF1WgyHy/Zt4G1h4UMCaSRHWO0jZJ/ayoJnQrr0C
lBQZL+LFMI3wlep+RKcWzCN2vpA8mGN3mQ9e+BNEwIxpaartrTyP57XCD4OnjEX9
G+/yTz2EWB5gNyPlPCiyHSTTuESHtttCxRG3TmxHWKSq70CpAPoSXKgW0uWAHMBp
bqihh7sF5ZIxm0jgquNzdPePJh5PpgjsFVTKoWgm3IQsvYEr9rn+7ccHGvRgiadu
FSUAbM1wxACBVlcKDwIFYVAaXrHL09OZthkw4gC+yK7k38km8lg/vsTlw7YucLm8
C4n+WkVA9PtDGJBGwZGshx20CP4iS8lE/LzrpYLhuEp0GT5fjoUvOuZRx9hfdWui
YRzIOsigerrfXfzIfzQ/6x1e2JwUe6aeRuSFhM8kpotXw9vseu9DYgoQgz8MOIjJ
gnSRnh/NNcAlyasfL/xs96D0rRQyGNotUL1B2quHLA83ZNk5nCZ4CdCcFOfrEi6h
kJu7M0KDJPsKaNBTPemiGcvMVtgeTAnYhrY1MZ1cHmsEgXmy2UkkYYJHcsyIZcsc
rzKax0etITI6ATFo45M1jJEZlHC3MEIqASkhXrs6pE+hUPbUBVCEFOJukUbmgTdI
lfT7Kn9Q+POug4Dn8J44fmB6MBA0DcROdL/VYHNm3yNS/G78/vYx6v5xHNrvb22E
KysPNMIY5V6LIw07mPk/2DzR5M+mbCew4fkE8X8PFuTBf96BH1E70Sq/F095JRgA
hrFqPmIWtGsdqJI94gyHZCZAwnDmnHjyWA+ARDMSQtwfVsig0LdWQdfRbWZMqGvP
QzfNul0jpvnFIWavcD6m+qG59uHkWwg0sUWezUr1fc5IS0Ou0xcuq/4L1ulrQmN4
aq6HHafCMZolJa0WQlhHHjTqoIkhYSbEefhqDz6N1JdlDpdCnZlLdtI80gvwL0h+
M9BOpFKLyuyWjweI6KJAagyYmQYzrI0tM1QqMhJc8GJ3DSM5wWrJTNGHUukshsbX
mTE6t6AVwnjAVY5ulRNrnR0QljzMlF67a74L3VYd3CRzFrVDSo3rtNoFHS1BA4nV
PJbx694faNvxlVTD9qQGynSP1KtSvBaAE2k2jUPPJl7gZLnr0HiNm8L8Jjyp1bml
BroLzsoBapNyoi+kJliDxbtboUwgkJE31VaV4YLqg6oljJWHtAOn83u4V9u5vlqi
Cn7H7v7sd1pOHTz69BYU4nebyBBcaBY3CpMeMq9KfFmXtoKEuorWQ7FiI31JAzZ7
j5A4bOGHsNPKrPB8DVr6rShYDwyK3PhIRLhWHRdWcGnk7eVTrcvwwSgsF8g8LGto
Y2ib1u5YO1sp2q3wPHW8CgVBq2XQk79mOCZKeTqlIY5eCnpTxmRrFyRo9eLahbgB
CE1Ezk/ZKzSMvEL5RStoiNGVWZPQNsbE1n6zbuuwDrpJ43gjlTXUkhb8aN/VUWwI
CO6Frhm1FlSjx4ueK/IA4SGiI7EFfHjnVm+vNhX1/BzTbDSXQ4M3B0g2KhieaBVi
4bULZbCH/flJXC1w/kgZirYsNDQM6j4Y7/EfVX6KPzywB5zlqnX0SpZN7mef420h
Hn7A8zzBa/YDSCxWNx2Gkq1USJ6ZA63Q0YDl/G9GFdE81P9gBYKJYgOiaVAOIo3G
4vTrSBWnrV1Ml6evJ9FxTFAOxcbRgYfG6RWG9xbKwUmTf/0jvs5Wpfc3ONv0cuhW
JLEkihqc3zIf+2Mu5GsJm/GPuBFvWqe56oyFuTqadkp6VbJsGn0bnbfC8ur6Txg5
Ld1fGb/cL2755I29BiVpJ1zRlFhNm71ipd5PsPRCACLBjtELbQrJRR5ewhYSGICA
/FUF59oN1hg5uFzUrcuJeRK/90xShlvYrPy35Yrnj8OUED19IDo62bArGl3/oSRc
3AgAsQ8qPtHyNyw0eZt3DyuJUdqmuz3+gqoEy4BoJkHz3/D6DjQs/3k2SMT9idBC
7PSrNw8GTkpAgmiPos2YkzIEh20myL+Kp/vqan7Diiuzc+cgYOT3JvhS+vRuUuMn
NYBNYsxCC0asR3TdvxjGROfrBk9k2+BFpdnof54BSP0IQCd+MfStRCw6fp/8oFMi
fYdrLZgdXbsiB6mhRvsHBd1uJd+Lpi63Wy8GTQ8Czdj2nyN/hkgNobPxJ3JelUD4
b2EaD6c2QLbMe8pNm5yJkWZiXA05SjUXSKp5CqV9ysrkFpt5NGDnItBrMUn6tcRX
Ll2MaFssjDbRUkay2C1o8o9aiEcc4rcobU19TCbk3/qPkvpMCLUDB0WO2Xp9ba+4
DgtiMT8CDjo306ScK9t5ps2BH3mLW9s41vX4WF/BiK21yZ3Z/nOnt+Fr/ky1AXfq
aYbHmVHQwiam7WnlD7IKBlOeUNtYgsQs9v2pe+XuBDNRCpKUWZd2y1tVJGoOFgHf
VU8QnLGRhcnwbFtfB9y/KsIep0iY3rf8Xawzz8jpqnCTlfSKOQQuo+aGTM2pSMZv
yMNX44K2xlisa4l7+G7NvAYMi3YBIvDHc3bf8uRFiLgg0dXUHGa0CsHm8269TBhD
n4DrGy9aN7ztfsJgRnxLmrv+dj7zKVDSBXNhy44af6NiXUI8H3PwgEv4L8d6R868
QmI8+YHPL6iZ0eYV/PgX+BO5X6yjPU3XfSGjp6ewuqIzeSAAq4wvC31rb1z6uRsv
iPFI59l5SLqD+IYkAQydqa+Jwr8hEbM72yarYXQKf7y41GBHZuUwTlcik7rLrZHs
eLXM6iqFSjm4GVABmZpANniSUpPmoO1wE/op8c9DMgVFX8mMvyH5kTeIwbHzVkzI
7ZGsGhA3Sp4qdpiPD01N6DDEupTD63DgR+iq+I+Ikr/r7ef6l975udpr95MmE2cU
FLBTqm4mKFPdVb0eBFaDJogl2IEbpyToRNuvOo9+yeAbrjDLkyU9NLHgXHptBMTd
4hbkQJSiRws6laSrYgZXUO5iWKAwFOHJJAhPVAfJdGis8BAAhi1YND9d1P0PL19O
ek77dI71AaN3w8EDJvwX4GBNKRQinKi2R+aCJkNOQCaHnH1or8s3Tv8Hr+TNxPFo
pV5GGQswKHYMuLt+nHMgqp/KOjv+FPLte2VQe/dQJ4F/YeGJIjziu0sfqaapWYOO
QcEwZiVr3SVYOFrPZ7ViXYYRW/8XUPgG1/7hZ74ovDyefLO4t4BiyO8tvJmhKtJq
h19vfKyAFMRRMzTFEIP5gxoT8DDweLcJa7rcWKgNYuMvHH0S/usgybh+4w3a/NHd
Q0PHAAzZ7hcLkrHWOLU8TnbkQzBg31Mje4T0MkDHKXtuESYYafhJHKQOVC7Tuip3
PZroTp6QG8iUFNUw8nFdXh1gky3sjieUgK3hNqXXYXoyt1KNdV+zZBHaARxbuoln
OQBPnu1lJShTxJ7PXnEwc8yrlZE1qkRjy9GTcd2KCo1Fn+RfX+Ehf9iDYwhyrsiX
/7G3ivuG16x5U7vTqwDwuAm+L88iQKrH2R2TtmRdZzJ1aJCOGE0REz+gCa4a7d6y
QMf67W3EYzeomf8zvHFxm5lTAGvhnzxAMuLuzHiQf23Tr9ahewcd77vCvh7qQJ6E
cgRUBaAx9Vbok9sOIvNEYjnXeHKVYdp8xAJXY7beyCq9XagGehZJ70VS4RALch67
QnQLJvLP+9nqgGXfkm73sLwLBg7i7kExGWytmm2S9hspjFqToWoRc8+zxGGRbNea
gmSFonp8xIoKPbQtK3QLSjPEFTo/kM4/smoaPvZ7F0ys0s885aj0lIae/hV67Hyn
y4PxYlz0Qv8wue9eV73jhgxN2L5dbKM2WLlKoFeTpTkXVeeWSwpDkKcJSzB50hDD
oU1zgOE35BlmJwjbv42UdfofQ2vE0k02psmBAdjbSj2PvogRFJGsAVyYzZumcrCS
/38YuQuc+vkdbmJDp+V+8t53kGIiD1s9KIEWFsOhLz3K67l7t1LcH2dkwfoPIcZA
Uexu9baSasLq1p+uGe8vAQeDmwE/cgNvSVGzOXq4rDv84rmb4ry7+HR8dgUdqXM5
TrqSIehXl4EpUSY7mzyOfNusIr0KbbqOCDbQD5GK1R400CD14xCv0TbuqxvnAbl1
RR5x3wUWHRm4v80dH+x8BDlAsbkffuzLIPoWk4dipxamJ1jmH1+fIpfI7ScXWg5C
mgN11asM1QcwLpx20HTPd34cD+2maz6uCWrLPkloXLQkD+rOtKsXsRw9Gk71XTmh
9K/NZp4R58eVAjBd5joJEhk5EDuL9Pj/uNW1erfXDPb9sSsnraVlOGQJuLUTHiqb
xMqplSf/tp/F48Qw0yjoXntPx5RX7RiUd+QlgJf3BLl+lqvKKasnfQaiQSPxKN/u
+EDU5cJi/4FIAk1WWtBnOm6UVZmfC+5gkEM5OfRLagvR/id5+zabz0uj5qQelBo/
xSbzWX+90VTsl7AxlhOmIZAhEqIiRB/pWkhHoUogZClUm1qvBfy7mpo2zQc2O6cA
jdO0K4OklLWmNhXCILUj8YtoDC5/apJqTx9AvdHvbTbNuwpGlXSqWKQ9mzrZv0Pp
E9G++MKJ0BRKAOQwJ/P9vfmtOrbyXdKqI4TF7Rtgtb6c8eX2kTrgRfK442SJtilC
etFXq8to5TbHcUlMllIYjX4P15dtRJEBN1UVYUjuxM/KT4eWnjcTf/JYbu5TO4Mt
/GS+lqcdNJb3pC0qT9ScEz1O0CP6OaypuKwtBeQryXs776WUeWCCTaiZC+Q5523J
ssfXCMRXCWjqj01DzUWjKsHxgCZm5bPGIUeNuZJrEemjPDI+fMourt0OLk6NULgg
rT4knkg+lo5E5EGNU2bIH+XV59XwhWYFA0gfkQY9+lIVaGVBuM8E5DcnpOvHYJb2
8UDT7QAmY7d457nHAxPoHz1fKR2JiMLbSbVoto+f6SWid/HNT/z3SXbd7dWB1Y2g
V3tZsiFseMlivlhegxZ7ZotyqlGsfjtk2ccm9quDaxuYRoQoA9uL1/QOpxdyBqWr
LISOP+nKa9y5xvCHKGIiOLatRy1bJWK8+ndRstiZ4PnHvzbH0nT8wpfd7rC4EB5I
scHHQ0cS6cvT8DlBNzn3yKSYYvjMHVhrLNp9pRWSpwAUu5kZ/hNcz33/NS8MpkK1
lTzHfMJrR++Gq8DOB0UD8/m8pX/Jr1eb1Ov5v0mQRCbS2ZckHzeaMaZbmuRhYQEN
1mb5EOIsOF91yNgpIgMYiuwf28XmiUn+6FIyABnjHovnxGPpCwJ818WWPqw46BGo
01rMXpfRQE7w0OjYmEerO2Hrl2K0Fp0M085tLg4+aFfzZ362fEsIZZPO2AA2kiMV
V8K/zcHoA+h9siTsbYVnSDAunxnXEHCIUYh7Su1XjAgS4aDHEJ8PWoMQv/mgtsls
N1jGvmg4SVJBxH7k9X+dcNaUaQ3OarQ5WrTOtNEUwkgEhHHSJcu3Kuc+19MaS8Am
L47LEnf/hbAi3HRPPgvzMjkbWkatElhWi4SirfLOBByjVkK2tlYfknKWtinfmTFw
SsnAQxvdXtrW+p4BqWX1F7+uzp9kP5V8WZy9RWe9U2QGUMRL/cFvL6LGE7rl7fac
FHhmpe78xOV5sN2NCvl7tnrii5zzxKWw1nrwd5wNwA6kaTPatO1VugVQTx5cQ6ia
Hp9rrLe5xv5ItOAzi2DO8Q6UX5CjDSMPjWKYF6OPr876Tqq9u8ZqjtahdhgfUfJe
aGycQ/NyogAJ/VQQLnivLf/c9XTll/QMXFve6wUwRmEMlPDtq0UsGvYyVuboUJr3
PGywfgWeJ3lPd+3hwcWHw3Pow0+eum1Bgpl2n/hr4CLIBQbbMpZ+M8sa8QX05dFS
ZXDOg6iL5HHKio8LAxy9VDqMbbg4JI/veIZivD7R8g5Y6Mm1LRJ2V1POho0hmlth
z/hq8Joz+zgYqO+o65bPqgN+MPJ1seFMoGIEKsBrTQVCpfX6rt7u459awdlIEysZ
EYVqKWaqRgLi2Ai18Cdc4hj3aqtoanbofksXfKaO+An9gzoSt+BoKvUXSXE9k7nc
3Qj1b9FcNoA+ZLXycmPDhTMpgZcmZftleF7pIxtw6Xkitqwrc1toZdJI/3gNANYU
lT15o87pxRHz8svXkOcyxmeAEx96Di6Q3P43b0HfCvmPU8nFNR7DUSuIsqMtcK6P
yVxDr80eR3BYO2tqGCKUFhsZqlsO5v7YcFCnMhhz/JEY8RoQZ2Kv2qokupPXukOm
3ahxnJgyHIP7wyBsFdgp24EOrA+O+R2Pkq54GERhHEU=
`pragma protect end_protected
